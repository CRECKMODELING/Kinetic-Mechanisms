   THERMO 
   300.0   1000.0   3000.0
CELL                    C   6H  10O   5     S 300.0    4000.0    1000.0        1
 2.92516210e+01 1.95010807e-02 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-1.25919988e+05 0.00000000e+00 2.92516210e+01 1.95010807e-02 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-1.25919988e+05 0.00000000e+00                   4
GMSW                    C   5H   8O   4     S 300.0    4000.0    1000.0        1
 2.38346742e+01 1.58897828e-02 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-1.03039895e+05 0.00000000e+00 2.38346742e+01 1.58897828e-02 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-1.03039895e+05 0.00000000e+00                   4
XYHW                    C   5H   8O   4     S 300.0    4000.0    1000.0        1
 2.38346742e+01 1.58897828e-02 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-1.07071125e+05 0.00000000e+00 2.38346742e+01 1.58897828e-02 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-1.07071125e+05 0.00000000e+00                   4
XYGR                    C   5H   8O   4     S 300.0    4000.0    1000.0        1
 2.38346742e+01 1.58897828e-02 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-1.09720219e+05 0.00000000e+00 2.38346742e+01 1.58897828e-02 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-1.09720219e+05 0.00000000e+00                   4
LIGC                    C  15H  14O   4     S 300.0    4000.0    1000.0        1
 4.65946547e+01 3.10631031e-02 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-1.03601488e+05 0.00000000e+00 4.65946547e+01 3.10631031e-02 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-1.03601488e+05 0.00000000e+00                   4
LIGH                    C  22H  28O   9     S 300.0    4000.0    1000.0        1
 7.87405700e+01 5.24937133e-02 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-2.24303494e+05 0.00000000e+00 7.87405700e+01 5.24937133e-02 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-2.24303494e+05 0.00000000e+00                   4
LIGO                    C  20H  22O  10     S 300.0    4000.0    1000.0        1
 7.62020414e+01 5.08013609e-02 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-2.51966073e+05 0.00000000e+00 7.62020414e+01 5.08013609e-02 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-2.51966073e+05 0.00000000e+00                   4
TGL                     C  57H 100O   7     S 300.0    4000.0    1000.0        1
 1.61902232e+02 1.07934821e-01 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-2.44625348e+05 0.00000000e+00 1.61902232e+02 1.07934821e-01 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-2.44625348e+05 0.00000000e+00                   4
TANN                    C  15H  12O   7     S 300.0    4000.0    1000.0        1
 5.48900197e+01 3.65933465e-02 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-1.59515809e+05 0.00000000e+00 5.48900197e+01 3.65933465e-02 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-1.59515809e+05 0.00000000e+00                   4
MOIST                   C   0H   2O   1     S 300.0    4000.0    1000.0        1   !From DH vaporization  engineering tool box
 9.04470000E+00 1.60000000E-03-6.00000000E-06 6.00000000E-09-2.00000000E-12    2
-3.70865499E+04-2.88280137E+02 9.04470000E+00 1.60000000E-03-6.00000000E-06    3
 6.00000000E-09-2.00000000E-12-3.70865499E+04-2.88280137E+02                   4
ASH                     C   0H   0K   1     S 300.0    4000.0    1000.0        1
 1.80625030E+01 1.20416687E-02 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
-1.55939610E+04 0.00000000E+00 1.80625030E+01 1.20416687E-02 0.00000000E+00    3
 0.00000000E+00	0.00000000E+00-1.55939610E+04 0.00000000E+00                   4
CELLA                   C   6H  10O   5     S 300.0    4000.0    1000.0        1
 2.92516210e+01 1.95010807e-02 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-1.25919988e+05 0.00000000e+00 2.92516210e+01 1.95010807e-02 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-1.25919988e+05 0.00000000e+00                   4
HCE1                    C   5H   8O   4     S 300.0    4000.0    1000.0        1
 2.38346742e+01 1.58897828e-02 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-9.92237373e+04 0.00000000e+00 2.38346742e+01 1.58897828e-02 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-9.92237373e+04 0.00000000e+00                   4
HCE2                    C   5H   8O   4     S 300.0    4000.0    1000.0        1
 2.38346742e+01 1.58897828e-02 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-1.10741538e+05 0.00000000e+00 2.38346742e+01 1.58897828e-02 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-1.10741538e+05 0.00000000e+00                   4
LIGCC                   C  15H  14O   4     S 300.0    4000.0    1000.0        1
 4.65946547e+01 3.10631031e-02 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-7.69910033e+04 0.00000000e+00 4.65946547e+01 3.10631031e-02 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-7.69910033e+04 0.00000000e+00                   4
LIGOH                   C  19H  22O   8     S 300.0    4000.0    1000.0        1
 6.82624420e+01 4.55082946e-02 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-1.86693370e+05 0.00000000e+00 6.82624420e+01 4.55082946e-02 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-1.86693370e+05 0.00000000e+00                   4
LIG                     C  11H  12O   4     S 300.0    4000.0    1000.0        1
 3.75634032e+01 2.50422688e-02 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-9.42255209e+04 0.00000000e+00 3.75634032e+01 2.50422688e-02 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-9.42255209e+04 0.00000000e+00                   4
ITANN                   C   8H   4O   4     S 300.0    4000.0    1000.0        1
 2.96079278e+01 1.97386186e-02 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-9.52526629e+04 0.00000000e+00 2.96079278e+01 1.97386186e-02 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-9.52526629e+04 0.00000000e+00                   4
CHAR                    C   1               S 300.0    4000.0    1000.0        1
-1.00796361E-01	4.99828606E-03 0.00000000E+00 0.00000000E+00 0.00000000E+00    2           
-1.94683964E+02 0.00000000E+00-1.00796361E-01 4.99828606E-03 0.00000000E+00    3
 0.00000000E+00	0.00000000E+00-1.94683964E+02 0.00000000E+00                   4 
CHARO                   C   1H   0O   1     S 300.0    4000.0    1000.0        1
-1.00796361E-01	4.99828606E-03 0.00000000E+00 0.00000000E+00 0.00000000E+00    2           
-1.94683964E+02 0.00000000E+00-1.00796361E-01 4.99828606E-03 0.00000000E+00    3
 0.00000000E+00	0.00000000E+00-1.94683964E+02 0.00000000E+00                   4 
COH2S                   C   1H   2O   1     S 300.0    4000.0    1000.0        1
 5.41694681e+00 3.61129787e-03 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-4.28130513e+04 0.00000000e+00 5.41694681e+00 3.61129787e-03 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-4.28130513e+04 0.00000000e+00                   4
CO2S                    C   1H   0O   2     S 300.0    4000.0    1000.0        1
 7.93959940e+00 5.29306627e-03 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-4.00155073e+04 0.00000000e+00 7.93959940e+00 5.29306627e-03 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-4.00155073e+04 0.00000000e+00                   4
COS                     C   1H   0O   1     S 300.0    4000.0    1000.0        1
 5.05324318e+00 3.36882879e-03 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-9.45019792e+03 0.00000000e+00 5.05324318e+00 3.36882879e-03 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-9.45019792e+03 0.00000000e+00                   4
COSTIFFS                C   1H   0O   1     S 300.0    4000.0    1000.0        1
 5.05324318e+00 3.36882879e-03 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-9.45019792e+03 0.00000000e+00 5.05324318e+00 3.36882879e-03 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-9.45019792e+03 0.00000000e+00                   4
CH3OHS                  C   1H   4O   1     S 300.0    4000.0    1000.0        1
 5.78065044e+00 3.85376696e-03 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-2.63330830e+04 0.00000000e+00 5.78065044e+00 3.85376696e-03 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-2.63330830e+04 0.00000000e+00                   4
CH4S                    C   1H   4O   0     S 300.0    4000.0    1000.0        1
 2.89429422e+00 1.92952948e-03 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-9.21591184e+03 0.00000000e+00 2.89429422e+00 1.92952948e-03 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-9.21591184e+03 0.00000000e+00                   4
C2H4S                   C   2H   4O   0     S 300.0    4000.0    1000.0        1
 5.06118118e+00 3.37412079e-03 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
 4.92120269e+03 0.00000000e+00 5.06118118e+00 3.37412079e-03 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00 4.92120269e+03 0.00000000e+00                   4
C6H5OHS                 C   6H   6O   1     S 300.0    4000.0    1000.0        1
 1.69787889e+01 1.13191926e-02 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-1.86144892e+04 0.00000000e+00 1.69787889e+01 1.13191926e-02 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-1.86144892e+04 0.00000000e+00                   4
CH2OS                   C   1H   2O   1     S 300.0    4000.0    1000.0        1
 5.41694681e+00 3.61129787e-03 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-2.45084187e+04 0.00000000e+00 5.41694681e+00 3.61129787e-03 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-2.45084187e+04 0.00000000e+00                   4
H2S                     C   0H   2O   0     S 300.0    4000.0    1000.0        1
 3.63703630e-01 2.42469087e-04 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
 1.09946128e+03 0.00000000e+00 3.63703630e-01 2.42469087e-04 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00 1.09946128e+03 0.00000000e+00                   4
C2H6S                   C   2H   6O   0     S 300.0    4000.0    1000.0        1
 5.42488481e+00 3.61658988e-03 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-1.10454007e+04 0.00000000e+00 5.42488481e+00 3.61658988e-03 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-1.10454007e+04 0.00000000e+00                   4
VANILLIN                C   8H   8O   3     G    300.00   3500.00 1260.00      1
 1.36544650e+01 4.84143232e-02-2.42641798e-05 5.50487829e-09-4.76001947e-13    2
-5.18855416e+04-3.54575728e+01-4.86637458e+00 1.07210639e-01-9.42597942e-05    3
 4.25395949e-08-7.82416000e-12-4.72182900e+04 5.81751551e+01                   4
CRESOL                  C   7H   8O   1     G    300.00   4000.00 1000.00      1
 .109411883E+02 .359221340E-01-.155859930E-04 .305336930E-08-.221926260E-12    2
-.211837368E+05-.322120090E+02-.410479790E+01 .823735850E-01-.680002460E-04    3
 .287114670E-07-.487123580E-11-.173767210E+05 .440872850E+02                   4
N2                G 8/02N   2    0    0    0G   200.000  6000.00  1000.00      1
 2.95257637E+00 1.39690040E-03-4.92631603E-07 7.86010195E-11-4.60755204E-15    2
-9.23948688E+02 5.87188762E+00 3.53100528E+00-1.23660988E-04-5.02999433E-07    3
 2.43530612E-09-1.40881235E-12-1.04697628E+03 2.96747038E+00 0.00000000E+00    4
O2                ATcT3EO   2    0    0    0G    200.00   6000.00 1000.00      1	
 3.65980488E+00 6.59877372E-04-1.44158172E-07 2.14656037E-11-1.36503784E-15    2
-1.21603048E+03 3.42074148E+00 3.78498258E+00-3.02002233E-03 9.92029171E-06    3
-9.77840434E-09 3.28877702E-12-1.06413589E+03 3.64780709E+00 0.00000000E+00    4
C2H6                    C   2H   6          G    300.00   4000.00 1000.00      1
 .404666411E+01 .153538802E-01-.547039485E-05 .877826544E-09-.523167531E-13    2
-.124473499E+05-.968698313E+00 .429142572E+01-.550154901E-02 .599438458E-04    3
-.708466469E-07 .268685836E-10-.115222056E+05 .266678994E+01                   4
C6H5OH                  C   6H   6O   1     G    300.00   4000.00 1000.00      1
 .141552427E+02 .199350340E-01-.718219540E-05 .116229002E-08-.697147483E-13    2
-.181287441E+05-.517984911E+02-.290978575E+00 .408562397E-01 .242829425E-04    3
-.714477617E-07 .346002146E-10-.134129780E+05 .268745637E+02                   4
C6H10O5                 C   6H  10O   5     G    300.00   4000.00 1000.00      1
 .279850422E+02 .264166682E-01-.913640739E-05 .142923991E-08-.833656585E-13    2
-.114313686E+06-.117754445E+03-.781241700E+01 .125424511E+00-.116271866E-03    3
 .544734561E-07-.100746170E-10-.103428291E+06 .690300863E+02                   4
C2H5OH     8/12/15      C   2H   6O   1    0G   300.000  5000.000 1402.000    21
 8.14483865E+00 1.28314052E-02-4.29052743E-06 6.55971721E-10-3.76506611E-14    2
-3.24005526E+04-1.86241126E+01 2.15805861E-01 2.95228396E-02-1.68271048E-05    3
 4.49484797E-09-4.02451543E-13-2.94851823E+04 2.45725052E+01                   4
C2H4                    C   2H   4          G    300.00   4000.00 1000.00      1
 .399182724E+01 .104833908E-01-.371721342E-05 .594628366E-09-.353630386E-13    2
 .426865851E+04-.269081762E+00 .395920063E+01-.757051373E-02 .570989993E-04    3
-.691588352E-07 .269884190E-10 .508977598E+04 .409730213E+01                   4
CH4               G 8/99C  1 H  4    0    0 G   200.000  6000.00  1000.00      1
 1.65326226E+00 1.00263099E-02-3.31661238E-06 5.36483138E-10-3.14696758E-14    2
-1.00095936E+04 9.90506283E+00 5.14911468E+00-1.36622009E-02 4.91453921E-05    3
-4.84246767E-08 1.66603441E-11-1.02465983E+04-4.63848842E+00-8.97226656E+03    4
C5H8O4                  C   5H   8O   4     G    300.00   4000.00 1000.00      1
 .217298154E+02 .217807665E-01-.749545594E-05 .116860895E-08-.680038942E-13    2
-.866505360E+05-.835752527E+02-.684199090E+01 .100610553E+00-.924172541E-04    3
 .429800586E-07-.789719358E-11-.779623201E+05 .655426910E+02                   4
HCOOH                   C   1H   2O   2     G    300.00   4000.00 1000.00      1   
 .461383160E+01 .644963640E-02-.229082510E-05 .367160470E-09-.218736750E-13    2
-.453303180E+05 .847883830E+00 .389836160E+01-.355877950E-02 .355205380E-04    3
-.438499590E-07 .171077690E-10-.467785744E+05 .734953970E+01                   4
CH3OH             T06/02C   1H  4 O  1    0 G   200.000  6000.00  1000.00      1
 3.52726795E+00 1.03178783E-02-3.62892944E-06 5.77448016E-10-3.42182632E-14    2
-2.60028834E+04 5.16758693E+00 5.65851051E+00-1.62983419E-02 6.91938156E-05    3
-7.58372926E-08 2.80427550E-11-2.56119736E+04-8.97330508E-01-2.41746056E+04    4
H2                ATcT3EH   2    0    0    0G    200.00   6000.00 1000.00      1
 2.90207649E+00 8.68992581E-04-1.65864430E-07 1.90851899E-11-9.31121789E-16    2
-7.97948726E+02-8.45591320E-01 2.37694204E+00 7.73916922E-03-1.88735073E-05    3
 1.95517114E-08-7.17095663E-12-9.21173081E+02 5.47184736E-01 0.00000000E+00    4
H2O               ATcT3EH   2O   1    0    0G    200.00   6000.00 1000.00      1
 2.73117512E+00 2.95136995E-03-8.35359785E-07 1.26088593E-10-8.40531676E-15    2
-2.99169082E+04 6.55183000E+00 4.20147551E+00-2.05583546E-03 6.56547207E-06    3
-5.52906960E-09 1.78282605E-12-3.02950066E+04-8.60610906E-01-2.90858262E+04    4
CO2               ATcT3EC   1O   2    0    0G    200.00   6000.00 1000.00      1
 4.63537470E+00 2.74559459E-03-9.98282389E-07 1.61013606E-10-9.22018642E-15    2
-4.90203677E+04-1.92887630E+00 2.20664321E+00 1.00970086E-02-9.96338809E-06    3
 5.47155623E-09-1.27733965E-12-4.83529864E+04 1.05261943E+01-4.73241678E+04    4
CO                ATcT3EC   1O   1    0    0G    200.00   6000.00 1000.00      1
 3.03397274E+00 1.37328118E-03-4.96445087E-07 8.10281447E-11-4.85331749E-15    2
-1.42586044E+04 6.10076092E+00 3.59508377E+00-7.21196937E-04 1.28238234E-06    3
 6.52429293E-10-8.21714806E-13-1.43448968E+04 3.44355598E+00-1.32928623E+04    4
CH2O                    C   1H   2O   1     G    300.00   4000.00 1000.00      1
 .316952665E+01 .619320560E-02-.225056366E-05 .365975660E-09-.220149458E-13    2
-.145486831E+05 .604207898E+01 .479372312E+01-.990833322E-02 .373219990E-04    3
-.379285237E-07 .131772641E-10-.143791953E+05 .602798058E+00                   4
C2H5CHO                 C   3H   6O   1     G    300.00   4000.00 1000.00      1
 .744085690E+01 .177301764E-01-.634081568E-05 .102040803E-08-.609461714E-13    2
-.260055814E+05-.144195446E+02 .424529681E+01 .668296706E-02 .493337933E-04    3
-.671986124E-07 .267262347E-10-.241473007E+05 .690738560E+01                   4
C6H6O3                  C   6H   6O   3     G    300.00   4000.00 1382.00      1
 .193892545E+02 .186134462E-01-.631148097E-05 .975462374E-09-.564561412E-13    2
-.492678935E+05-.716786498E+02 .598814621E+00 .618493802E-01-.438009436E-04    3
 .155531333E-07-.220506530E-11-.427313109E+05 .293828012E+02                   4
CH3CHO            L 8/88C  2 H  4 O   1   0 G   200.000  6000.00  1000.00      1
 0.54041108E+01 0.11723059E-01-0.42263137E-05 0.68372451E-09-0.40984863E-13    2
-0.22593122E+05-0.34807917E+01 0.47294595E+01-0.31932858E-02 0.47534921E-04    3
-0.57458611E-07 0.21931112E-10-0.21572878E+05 0.41030159E+01-0.19987949E+05    4
CH2OHCH2CHO             C   3H   6O   2     G    300.00   4000.00 1382.00      1
 .118936666E+02 .144153203E-01-.477525443E-05 .726036430E-09-.415285995E-13    2
-.459271652E+05-.327285750E+02 .266613285E+01 .346302298E-01-.214380719E-04    3
 .690469334E-08-.916939105E-12-.425706030E+05 .173358364E+02                   4
FURFURAL                C   5H   4O   2     G    300.00   4000.00 1000.00      1
 .159553578E+02 .122096134E-01-.419491662E-05 .654219009E-09-.381060338E-13    2
-.255664634E+05-.596830465E+02-.186260023E+01 .570946426E-01-.476338594E-04    3
 .197949337E-07-.326585828E-11-.197873020E+05 .347179869E+02                   4
CH3CO2H                 C   2H   4O   2     G    300.00   4000.00 1000.00      1
 .767084601E+01 .135152602E-01-.525874333E-05 .893184479E-09-.553180543E-13    2
-.557560970E+05-.154677315E+02 .278950201E+01 .999941719E-02 .342572245E-04    3
-.509031329E-07 .206222185E-10-.534752488E+05 .141053123E+02                   4
C24H28O4                C  24H  28O   4     G    300.00   4000.00 1398.00      1
 .495886732E+02 .844753396E-02 .385179844E-05-.232491508E-08 .315199759E-12    2
-.164047630E+05-.193448260E+03 .542487420E+01 .999122905E-01-.513976516E-04    3
-.430175388E-08 .876106788E-11-.572347637E+04 .356171545E+02                   4
C2H3CHO           KPS12 C   3H   4O   1    0G   300.000  5000.000 1398.000    01
 9.99155394E+00 9.82348001E-03-3.31203088E-06 5.09524422E-10-2.93821890E-14    2
-1.25303509E+04-2.85168883E+01 7.33844455E-01 3.17482671E-02-2.29599468E-05    3
 8.42104232E-09-1.23613478E-12-9.38473548E+03 2.10308851E+01                   4
C6H5OCH3                C   7H   8O   1     G    300.00   4000.00 1393.00      1
 .203938728E+02 .209088165E-01-.722522263E-05 .112997840E-08-.659097524E-13    2
-.186061425E+05-.862920505E+02-.540888697E+01 .873332441E-01-.739639658E-04    3
 .320208039E-07-.556946955E-11-.102821510E+05 .500696056E+02                   4
U2ME12                  C  13H  22O   2     G    300.00   4000.00 1391.00      1
 .422353117E+02 .524987045E-01-.181261023E-04 .283174793E-08-.165001495E-12    2
-.676968189E+05-.186270028E+03 .679798314E-01 .152530074E+00-.111376081E-03    3
 .435663556E-07-.715842617E-11-.529996239E+05 .399987338E+02                   4
MLINO                   C  19H  34O   2     G    300.00   4000.00 1833.00      1
 .524257963E+02 .910351615E-01-.326514183E-04 .524998946E-08-.312507814E-12    2
-.869039436E+05-.227879204E+03-.158761924E+01 .219526542E+00-.145761172E-03    3
 .495347572E-07-.688636525E-11-.693288124E+05 .600962817E+02                   4
CH2OHCHO                C   2H   4O   2     G    300.00   4000.00 1000.00      1
 .691088832E+01 .123280849E-01-.438373062E-05 .703055164E-09-.419009846E-13    2
-.400211587E+05-.696132551E+01 .614926095E+01-.596828114E-02 .596003337E-04    3
-.716663578E-07 .274014411E-10-.388356849E+05 .186644598E+01                   4
CHOCHO                  C   2H   2O   2     G    300.00   4000.00 1000.00      1
 .872506895E+01 .633096819E-02-.235574814E-05 .389782853E-09-.237486912E-13    2
-.291024131E+05-.203903909E+02 .468412461E+01 .478012819E-03 .426390768E-04    3
-.579018239E-07 .231669328E-10-.271985007E+05 .451187184E+01                   4
HOCHO                   H   2C   1O   2     G    200.00   3500.00 1800.00      1
 3.79473623e+00 8.42765802e-03-3.84722303e-06 8.63389995e-10-7.73674578e-14    2
-4.73118220e+04 5.12934093e+00 1.85206267e+00 1.27447104e-02-7.44476667e-06    3
 2.19581357e-09-2.62426287e-13-4.66124595e+04 1.56434955e+01                   4
	
			     		  



