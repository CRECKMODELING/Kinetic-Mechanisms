! 
!
! A. Stagni, S. Arunthanayothin, L. Pratali Maffei,
! O. Herbinet, F. Battin-Leclerc, T. Faravelli
! "An experimental, theoretical and kinetic-modeling study of hydrogen sulfide pyrolysis and oxidation"
! Chemical Engineering Journal (submitted) (2022).
!
! Submitted to Chemical Engineering Journal (December 2021)
!
! Thermodynamic properties
! 
! CHEMKIN format
!
!VERSION:  17_03
!AUTHORS:  C1-C3   Burcat   
!NOTE:     SPECIES RE-ARRANGED AS THE SAME ORDER IN MECH
!
!VERSION:  17_05
!Following species are updated from ATcT's Database:
! H	H2	O	O2	HE
! OH	H2O	N2	HO2	HCO
! H2O2	AR	CO	CO2
 THERMO
  300.   1000.   4000.
HE                ATcT3EHe  1    0    0    0G    200.00   6000.00 1000.00      1 ! [Ghobad] He <g> ATcT ver. 1.122, DHf298 = 0.000 \B1 0.000 kJ/mol - fit MAR17
 2.49985609E+00 2.19365392E-07-1.07525085E-10 2.07198041E-14-1.39358612E-18    2
-7.45309155E+02 9.29535014E-01 2.49976293E+00 1.01013432E-06-8.24578465E-10    3
-6.85983306E-13 7.24751856E-16-7.45340917E+02 9.29800315E-01 0.00000000E+00    4
AR                ATcT3EAr  1    0    0    0G    200.00   6000.00 1000.00      1 ! [Ghobad] Ar <g> ATcT ver. 1.122, DHf298 = 0.000 \B1 0.000 kJ/mol - fit MAR17
 2.49989176E+00 1.56134837E-07-7.76108557E-11 1.52928085E-14-1.05304493E-18    2
-7.45328403E+02 4.38029835E+00 2.49988611E+00 2.13037960E-07 8.97320772E-10    3
-2.31395752E-12 1.30201393E-15-7.45354481E+02 4.38024367E+00 0.00000000E+00    4
N2                ATcT3EN   2    0    0    0G    200.00   6000.00 1000.00      1 ! [Ghobad] N2 <g> ATcT ver. 1.122, DHf298 = 0.000 \B1 0.000 kJ/mol - fit MAR17
 2.93802970E+00 1.41838030E-03-5.03281045E-07 8.07555464E-11-4.76064275E-15    2
-9.17180990E+02 5.95521985E+00 3.53603521E+00-1.58270944E-04-4.26984251E-07    3
 2.37542590E-09-1.39708206E-12-1.04749645E+03 2.94603724E+00 0.00000000E+00    4
O2                ATcT3EO   2    0    0    0G    200.00   6000.00 1000.00      1 ! [Ghobad] O2 <g> ATcT ver. 1.122, DHf298 = 0.000 \B1 0.000 kJ/mol - fit MAR17
 3.65980488E+00 6.59877372E-04-1.44158172E-07 2.14656037E-11-1.36503784E-15    2
-1.21603048E+03 3.42074148E+00 3.78498258E+00-3.02002233E-03 9.92029171E-06    3
-9.77840434E-09 3.28877702E-12-1.06413589E+03 3.64780709E+00 0.00000000E+00    4
H2                ATcT3EH   2    0    0    0G    200.00   6000.00 1000.00      1 ! [Ghobad] H2 <g> ATcT ver. 1.122, DHf298 = 0.000 \B1 0.000 kJ/mol - fit MAR17
 2.90207649E+00 8.68992581E-04-1.65864430E-07 1.90851899E-11-9.31121789E-16    2
-7.97948726E+02-8.45591320E-01 2.37694204E+00 7.73916922E-03-1.88735073E-05    3
 1.95517114E-08-7.17095663E-12-9.21173081E+02 5.47184736E-01 0.00000000E+00    4
H2O               ATcT3EH   2O   1    0    0G    200.00   6000.00 1000.00      1 ! [Ghobad] H2O <g> ATcT ver. 1.122, DHf298 = -241.833 \B1 0.027 kJ/mol - fit MAR17
 2.73117512E+00 2.95136995E-03-8.35359785E-07 1.26088593E-10-8.40531676E-15    2
-2.99169082E+04 6.55183000E+00 4.20147551E+00-2.05583546E-03 6.56547207E-06    3
-5.52906960E-09 1.78282605E-12-3.02950066E+04-8.60610906E-01-2.90858262E+04    4
H2O2              ATcT3EH   2O   2    0    0G    200.00   6000.00 1000.00      1 ! [Ghobad] H2O2 <g> ATcT ver. 1.122, DHf298 = -135.457 \B1 0.064 kJ/mol - fit MAR17
 4.54017480E+00 4.15970971E-03-1.30876777E-06 2.00823615E-10-1.15509243E-14    2
-1.79514029E+04 8.55881745E-01 4.23854160E+00-2.49610911E-04 1.59857901E-05    3
-2.06919945E-08 8.29766320E-12-1.76486003E+04 3.58850097E+00-1.62917334E+04    4
O                 ATcT3EO   1    0    0    0G    200.00   6000.00 1000.00      1 ! [Ghobad] O <g> ATcT ver. 1.122, DHf298 = 249.229 \B1 0.002 kJ/mol - fit MAR17
 2.55160087E+00-3.83085457E-05 8.43197478E-10 4.01267136E-12-4.17476574E-16    2
 2.92287628E+04 4.87617014E+00 3.15906526E+00-3.21509999E-03 6.49255543E-06    3
-5.98755115E-09 2.06876117E-12 2.91298453E+04 2.09078344E+00 2.99753606E+04    4
H                 ATcT3EH   1    0    0    0G    200.00   6000.00 1000.00      1 ! [Ghobad] H <g> ATcT ver. 1.122, DHf298 = 217.998 \B1 0.000 kJ/mol - fit MAR17
 2.49985211E+00 2.34582548E-07-1.16171641E-10 2.25708298E-14-1.52992005E-18    2
 2.54738024E+04-4.45864645E-01 2.49975925E+00 6.73824499E-07 1.11807261E-09    3
-3.70192126E-12 2.14233822E-15 2.54737665E+04-4.45574009E-01 2.62191345E+04    4
OH                ATcT3EH   1O   1    0    0G    200.00   6000.00 1000.00      1 ! [Ghobad] OH <g> ATcT ver. 1.122, DHf298 = 37.490 \B1 0.027 kJ/mol - fit MAR17
 2.84581721E+00 1.09723818E-03-2.89121101E-07 4.09099910E-11-2.31382258E-15    2
 3.71706610E+03 5.80339915E+00 3.97585165E+00-2.28555291E-03 4.33442882E-06    3
-3.59926640E-09 1.26706930E-12 3.39341137E+03-3.55397262E-02 4.50901087E+03    4
HO2               ATcT3EH   1O   2    0    0G    200.00   6000.00 1000.00      1 ! [Ghobad] HO2 <g> ATcT ver. 1.122, DHf298 = 12.26 \B1 0.16 kJ/mol - fit MAR17 
 4.10564010E+00 2.04046836E-03-3.65877562E-07 1.85973044E-11 4.98818315E-16    2
 4.32898769E+01 3.30808126E+00 4.26251250E+00-4.45642032E-03 2.05164934E-05    3
-2.35794011E-08 9.05614257E-12 2.62442356E+02 3.88223684E+00 1.47417835E+03    4
!+++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
!SOx MODULE
!+++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
S                 J 9/82S  1.   0.   0.   0.G   200.000  6000.000 1000.        1 ! Burcat database http://garfield.chem.elte.hu/Burcat/THERM.DAT
 2.87936498E+00-5.11050388E-04 2.53806719E-07-4.45455458E-11 2.66717362E-15    2
 3.25013791E+04 3.98140647E+00 2.31725616E+00 4.78018342E-03-1.42082674E-05    3
 1.56569538E-08-5.96588299E-12 3.25068976E+04 6.06242434E+00 3.33128471E+04    4
S2                tpis89S  2.   0.   0.   0.G   200.000  6000.000 1000.        1 ! Burcat database http://garfield.chem.elte.hu/Burcat/THERM.DAT
 3.83249656E+00 8.88970881E-04-2.59080844E-07 3.63847115E-11-1.72606371E-15    2
 1.42836134E+04 5.33000845E+00 2.87736627E+00 5.00301430E-03-6.04370732E-06    3
 3.04738962E-09-3.87017618E-13 1.44342379E+04 9.79873919E+00 1.54669367E+04    4
SO                tpis89S  1.O  1.   0.   0.G   200.000  6000.000 1000.        1 ! Burcat database http://garfield.chem.elte.hu/Burcat/THERM.DAT
 3.96894225E+00 3.77296831E-04 7.67102696E-09-1.37544433E-11 1.37139416E-15    2
-7.28571725E+02 3.73493087E+00 3.61859514E+00-2.32173768E-03 1.16462669E-05    3
-1.42092510E-08 5.60765370E-12-4.80621641E+02 6.36504115E+00 5.72529951E+02    4
S2O               tpis89S  2.O  1.   0.   0.G   200.000  6000.000 1000.        1 ! Burcat database http://garfield.chem.elte.hu/Burcat/THERM.DAT
 6.02401811E+00 1.00035579E-03-3.91923038E-07 6.69240060E-11-4.16275707E-15    2
-8.76531218E+03-2.93690271E+00 3.01869800E+00 1.08575811E-02-1.25419070E-05    3
 6.57657832E-09-1.21573834E-12-8.02370855E+03 1.21738889E+01-6.73948254E+03    4
SO2               tpis89S  1.O  2.   0.   0.G   200.000  6000.000 1000.        1 ! Burcat database http://garfield.chem.elte.hu/Burcat/THERM.DAT
 5.38423482E+00 1.67930560E-03-6.32062944E-07 1.08465348E-10-6.66890336E-15    2
-3.76067022E+04-1.83130517E+00 3.67480752E+00 2.28302107E-03 8.46893049E-06    3
-1.36562039E-08 5.76271873E-12-3.69455073E+04 7.96866430E+00-3.56978343E+04    4
SO3               tpis89S  1.O  3.   0.   0.G   200.000  6000.000 1000.        1 ! Burcat database http://garfield.chem.elte.hu/Burcat/THERM.DAT
 7.29677572E+00 2.73576437E-03-1.06377755E-06 1.80776031E-10-1.12077527E-14    2
-5.03096739E+04-1.24246659E+01 2.37461122E+00 1.59543297E-02-1.26322543E-05    3
 2.81827264E-09 6.23371547E-13-4.89269231E+04 1.31043046E+01-4.76155540E+04    4
SH                IU2/03S  1.H  1.   0.   0.G   200.000  6000.000 1000.        1 ! Burcat database http://garfield.chem.elte.hu/Burcat/THERM.DAT
 3.03153027E+00 1.25805252E-03-4.05524133E-07 6.19648110E-11-3.50862111E-15    2
 1.62059674E+04 6.15022140E+00 3.68466877E+00 3.24608824E-03-1.28635079E-05    3
 1.69512196E-08-7.07595387E-12 1.59036477E+04 2.01781634E+00 1.70629418E+04    4
HS2 anharmonic    T 3/03H  1.S  2.   0.   0.G   200.000  6000.000 1000.        1 ! Burcat database http://garfield.chem.elte.hu/Burcat/THERM.DAT
 4.75155728E+00 2.15521745E-03-7.39343908E-07 1.22229939E-10-7.35968292E-15    2
 1.08214337E+04 2.68990027E+00 2.96279116E+00 8.56185025E-03-9.91987786E-06    3
 6.19874244E-09-1.52120491E-12 1.12507023E+04 1.15828502E+01 1.24384961E+04    4
HOS                SDT18 S  1 H  1 O  1     G    200.00   3000.00 1000.00      1 ! Fit from Glarborg et al. Int Jour Chem Kinet 28 (1996)
+3.70066631E+00+3.91895206E-03-2.62851749E-06+9.32360519E-10-1.19646656E-13    2
-1.29963559E+03+6.50634821E+00+3.34253914E+00+3.22329148E-03+2.51066588E-06    3
-5.82651580E-09+2.55383405E-12-1.15171631E+03+8.69086055E+00                   4
HSO  HS=O         T04/07H  1.S  1.O  1.   0.G   200.000  6000.000 1000.        1  ! Burcat database
 4.34724125E+00 2.53372236E-03-9.51430950E-07 1.58095446E-10-9.65294637E-15    2
-4.20893834E+03 3.15887502E+00 4.13565093E+00-3.69243127E-03 2.05169784E-05    3
-2.40530656E-08 9.17084270E-12-3.82371653E+03 5.88770120E+00-2.61672666E+03    4
HSO2               SDT18 S  1 H  1 O  2     G    200.00   3000.00 1000.00      1 ! Fit from Glarborg et al. Int Jour Chem Kinet 28 (1996)
+4.15733956E+00+1.04743749E-02-8.00819825E-06+2.82571970E-09-3.62209570E-13    2
-1.87567868E+04+5.31642597E+00+3.42869741E+00+8.42027402E-03+4.55829457E-06    3
-1.32303946E-08+5.91015498E-12-1.84303695E+04+9.90450909E+00                   4
HSOO               SDT18 H  1 S  1 O  2     G    298.00   3000.00 1000.00      1 ! Fit from Song et al. Int. J. Chem. Kinet. 49 37-52 (2017)
+4.41364109E+00+8.27319630E-03-6.12760846E-06+2.16146744E-09-2.76958440E-13    2
+1.46172646E+04+6.65022426E+00+3.81424283E+00+1.04127009E-02-8.18175865E-06    3
+2.24884699E-09+1.49705835E-13+1.47244496E+04+9.54249866E+00                   4
HOSO               SDT18 S  1 H  1 O  2     G    200.00   3000.00 1000.00      1 ! Fit from Glarborg et al. Int Jour Chem Kinet 28 (1996)
+5.21864278E+00+6.61085720E-03-4.68100796E-06+1.65149640E-09-2.11637427E-13    2
-3.09869415E+04+6.89488722E-01+3.56075878E+00+8.39294787E-03+2.05454098E-06    3
-1.05343375E-08+5.11444086E-12-3.04840430E+04+9.72230559E+00                   4
HOSO2              SDT18 S  1 H  1 O  3     G    200.00   3000.00 1000.00      1 ! Fit from Glarborg et al. Int Jour Chem Kinet 28 (1996)
+7.81496344E+00+7.40652535E-03-5.30611412E-06+1.87201113E-09-2.39895582E-13    2
-4.98551261E+04-1.13522005E+01+5.23391459E+00+1.16161683E-02+5.83624122E-07    3
-1.22121987E-08+6.32598193E-12-4.91342678E+04+2.37580849E+00                   4
H2S                     H   2S   1          G    300.00   5000.00 1000.00      1 ! Burcat database http://garfield.chem.elte.hu/Burcat/THERM.DAT
 .288314700E+01 .382783500E-02-.142339800E-05 .249799900E-09-.166027300E-13    2
-.348074300E+04 .725816200E+01 .307102900E+01 .557826100E-02-.103096700E-04    3
 .120195300E-07-.483837000E-11-.355982600E+04 .593522600E+01                   4
H2S2  H-S-S-H     T 3/03H  2.S  2.   0.   0.G   200.000  6000.000 1000.        1 ! Burcat database http://garfield.chem.elte.hu/Burcat/THERM.DAT
 5.69402902E+00 3.90495326E-03-1.41886468E-06 2.30688658E-10-1.38745854E-14    2
-1.65807167E+02-3.74138641E+00 2.09117166E+00 1.94220358E-02-2.89395611E-05    3
 2.30251562E-08-7.20187083E-12 5.91056782E+02 1.35883795E+01 1.86421088E+03    4
HSOH               SDT18 S  1 H  2 O  1     G    200.00   3000.00 1000.00      1 ! Fit from Glarborg et al. Int Jour Chem Kinet 28 (1996)
+3.22369152E+00+1.09195807E-02-8.34107303E-06+2.94324835E-09-3.77281906E-13    2
-1.58051933E+04+8.05599967E+00+3.54299277E+00+4.88607922E-03+9.18329891E-06    3
-1.52821960E-08+6.03799076E-12-1.56758945E+04+7.59299028E+00                   4
H2SO               SDT18 S  1 H  2 O  1     G    200.00   3000.00 1000.00      1 ! Fit from Glarborg et al. Int Jour Chem Kinet 28 (1996)
+7.28881818E-01+1.66806861E-02-1.27837855E-05+4.51059240E-09-5.78163226E-13    2
-6.54928648E+03+2.02124212E+01+2.67153709E+00+4.94767340E-03+1.19552752E-05    3
-1.75391118E-08+6.52283778E-12-6.77956309E+03+1.17311676E+01                   4
HOSHO              SDT18 S  1 H  2 O  2     G    200.00   3000.00 1000.00      1 ! Fit from Glarborg et al. Int Jour Chem Kinet 28 (1996)
+4.56801477E+00+1.32625658E-02-9.79156366E-06+3.45461897E-09-4.42738075E-13    2
-3.44927587E+04+2.50254289E+00+3.49309948E+00+1.04449987E-02+7.89362227E-06    3
-1.91633903E-08+8.38256771E-12-3.40146806E+04+9.23577879E+00                   4
END
