!"A comprehensive kinetic framework for solid carbon deposition and hydrogen production from the pyrolysis of light
!                                             hydrocarbons streams."
!                                        
!Francesco Serse (a), Zhaobin Ding �(b), Mauro Bracconi (b), Matteo Maestri �(b), Andrea Nobili (a), Clarissa Giudici (a), Alessio Frassoldati (a), Tiziano Faravelli (a),
!                                       Alberto Cuoci (a), Matteo Pelucchi* (a).
!                                        
!               a) CRECK Modelling Lab, Department of Chemistry Materials and Chemical Engineering, Politecnico di Milano, Italy.
!               b) LCCP Department of Energy, Politecnico di Milano, Italy.
!               � current affiliation: School of Chemical Engineering and Technology, Sun Yat-Sen University (SYSU), Guangzhou, China.


                                        
!Corresponding authors:
!*matteo.pelucchi@polimi.it
!�matteo.maestri@polimi.it


! This thermodynamic database was obtained by fitting the thermodynamic properties
! extracted from the following file: TOT2003.THERM
! The thermodynamic properties are fitted in order to preserve not only the 
! continuity of each function at the intermediate temperature, but also the  continuity
! of the derivatives, from the 1st to the 3rd order
! The intermediate temperatures are chosen in order to minimize the fitting error.
! Last update: 3/25/2020

THERMO ALL
270.   1000.   3500. 
AR                      AR  1               G    200.00   3500.00  820.00      1
 2.50013931e+00-3.98290200e-07 3.45886082e-10-1.18293971e-13 1.38553174e-17    2
-7.45407891e+02 4.37897362e+00 2.49974489e+00 1.52569132e-06-3.17359231e-09    3
 2.74307057e-12-8.58511922e-16-7.45343207e+02 4.38079817e+00                   4
N2                      N   2               G    200.00   3500.00 1050.00      1
 2.81166073e+00 1.67067353e-03-6.79997428e-07 1.32881379e-10-1.02767442e-14    2
-8.69811579e+02 6.64838050e+00 3.73100682e+00-1.83159730e-03 4.32324662e-06    3
-3.04378151e-09 7.46071562e-13-1.06287426e+03 2.16821198e+00                   4
HE                      HE  1               G    200.00   3500.00  850.00      1
 2.50020615e+00-5.42576298e-07 4.63926302e-10-1.57302170e-13 1.82971406e-17    2
-7.45426807e+02 9.27648988e-01 2.49964853e+00 2.08151569e-06-4.16682427e-09    3
 3.47465907e-12-1.04992675e-15-7.45332012e+02 9.30248556e-01                   4
H2                      H   2               G    200.00   3500.00  700.00      1
 3.78199881e+00-1.01873259e-03 1.24226233e-06-4.19011898e-10 4.75543793e-14    2
-1.10283023e+03-5.60525910e+00 2.64204438e+00 5.49529274e-03-1.27163634e-05    3
 1.28749173e-08-4.70027749e-12-9.43236614e+02-5.12231102e-01                   4
H                       H   1               G    200.00   3500.00  860.00      1
 2.50031493e+00-7.73406828e-07 6.39345346e-10-2.12551791e-13 2.44479191e-17    2
 2.54736474e+04-4.48357228e-01 2.49950544e+00 2.99164046e-06-5.92759759e-09    3
 4.87810165e-12-1.45539320e-15 2.54737866e+04-4.44574018e-01                   4
O2                      O   2               G    200.00   3500.00  700.00      1
 2.82012408e+00 2.48211357e-03-1.51202094e-06 4.48556201e-10-4.87305668e-14    2
-9.31350148e+02 7.94914552e+00 3.74403921e+00-2.79740147e-03 9.80122558e-06    3
-1.03259643e-08 3.79931247e-12-1.06069827e+03 3.82132646e+00                   4
O                       O   1               G    200.00   3500.00  720.00      1
 2.62549143e+00-2.08959644e-04 1.33918546e-07-3.85875896e-11 4.38918689e-15    2
 2.92061519e+04 4.48358519e+00 3.14799201e+00-3.11174065e-03 6.18137897e-06    3
-5.63808798e-09 1.94866016e-12 2.91309118e+04 2.13446549e+00                   4
H2O                     H   2O   1          G    200.00   3500.00 1420.00      1
 2.66777075e+00 3.05768849e-03-9.00442411e-07 1.43361552e-10-1.00857817e-14    2
-2.98875645e+04 6.91191131e+00 4.06061172e+00-8.65807189e-04 3.24409528e-06    3
-1.80243079e-09 3.32483293e-13-3.02831314e+04-2.96150481e-01                   4
OH                      H   1O   1          G    200.00   3500.00 1700.00      1
 2.49867369e+00 1.66635279e-03-6.28251516e-07 1.28346806e-10-1.05735894e-14    2
 3.88110716e+03 7.78218862e+00 3.91354631e+00-1.66275926e-03 2.30920029e-06    3
-1.02359508e-09 1.58829629e-13 3.40005047e+03 2.05474719e-01                   4
H2O2                    H   2O   2          G    200.00   3500.00 1800.00      1
 4.76869639e+00 3.89237848e-03-1.21382349e-06 1.92615285e-10-1.22581990e-14    2
-1.80900220e+04-5.11811777e-01 3.34774224e+00 7.05005437e-03-3.84522006e-06    3
 1.16720661e-09-1.47618105e-13-1.75784785e+04 7.17868851e+00                   4
HO2                     H   1O   2          G    200.00   3500.00  700.00      1
 3.02391889e+00 4.46390907e-03-2.23146492e-06 6.12710799e-10-6.64266237e-14    2
 3.99341609e+02 9.10699973e+00 3.61994299e+00 1.05805705e-03 5.06678941e-06    3
-6.33800762e-09 2.41597281e-12 3.15898234e+02 6.44411482e+00                   4
CO                      C   1O   1          G    200.00   3500.00  960.00      1
 2.79255381e+00 1.87486886e-03-8.59711926e-07 1.91200070e-10-1.67855286e-14    2
-1.41723335e+04 7.41443560e+00 3.75723891e+00-2.14465241e-03 5.42079005e-06    3
-4.17025963e-09 1.11901127e-12-1.43575530e+04 2.79976799e+00                   4
CO2                     C   1O   2          G    200.00   3500.00 1450.00      1
 4.70876468e+00 2.62914704e-03-9.30606462e-07 1.43892920e-10-7.62581414e-15    2
-4.90562639e+04-2.34976452e+00 2.31684347e+00 9.22755036e-03-7.75654093e-06    3
 3.28225360e-09-5.48722482e-13-4.83626067e+04 1.00786234e+01                   4
HOCO                    H   1C   1O   2     G    200.00   3500.00 1570.00      1
 5.88810541e+00 3.28985507e-03-9.88703861e-07 1.12295277e-10-2.32818718e-15    2
-2.40914384e+04-5.05613727e+00 2.36661498e+00 1.22618052e-02-9.56063074e-06    3
 3.75217930e-09-5.81927554e-13-2.29856904e+04 1.35214769e+01                   4
CH4                     C   1H   4          G    300.00   3500.00  700.00      1
 5.05346405e-01 1.23697845e-02-4.99807922e-06 1.04392765e-09-8.62897416e-14    2
-9.58982501e+03 1.61752775e+01 5.23967335e+00-1.46835123e-02 5.29732711e-05    3
-5.41668822e-08 1.96318566e-11-1.02526308e+04-4.97649748e+00                   4
CH3                     C   1H   3          G    300.00   3500.00 1060.00      1
 2.78805104e+00 6.15233477e-03-2.21179349e-06 3.74402648e-10-2.48151349e-14    2
 1.65862829e+04 5.77899818e+00 3.47829310e+00 3.54764773e-03 1.47408440e-06    3
-1.94375955e-09 5.21921232e-13 1.64399516e+04 2.40875956e+00                   4
CH2                     C   1H   2          G    300.00   3500.00 1800.00      1
 2.81272972e+00 3.55431388e-03-1.28768523e-06 2.21273744e-10-1.48738147e-14    2
 4.62073492e+04 6.64284652e+00 3.76489460e+00 1.43839191e-03 4.75583077e-07    3
-4.31788591e-10 7.58292874e-14 4.58645699e+04 1.48953153e+00                   4
CH2(S)                  C   1H   2          G    300.00   3500.00  970.00      1
 2.75934299e+00 3.65468307e-03-1.35589914e-06 2.74980411e-10-2.36795472e-14    2
 5.06429079e+04 6.11646383e+00 4.18185434e+00-2.21134314e-03 7.71527541e-06    3
-5.95950381e-09 1.58314628e-12 5.03669407e+04-7.03002602e-01                   4
C                       C   1               G    200.00   3500.00  700.00      1
 2.49472531e+00 3.92839476e-05-6.70014980e-08 3.71818694e-11-5.07306885e-15    2
 8.54504422e+04 4.79314254e+00 2.54495192e+00-2.47725281e-04 5.48018277e-07    3
-5.48551250e-10 2.04117331e-13 8.54434105e+04 4.56874273e+00                   4
CH                      C   1H   1          G    300.00   3500.00 1590.00      1
 2.27990128e+00 2.16985238e-03-7.07637885e-07 1.23973494e-10-9.56348515e-15    2
 7.11059412e+04 8.77326061e+00 3.77264332e+00-1.58547350e-03 2.83512238e-06    3
-1.36146058e-09 2.23995332e-13 7.06312492e+04 8.79407904e-01                   4
CH3O2H                  C   1H   4O   2     G    300.00   3500.00 1090.00      1
 7.33435519e+00 9.33238534e-03-3.40995713e-06 5.79327692e-10-3.79241109e-14    2
-1.81046374e+04-1.19553974e+01 7.70006797e-01 3.34217373e-02-3.65604414e-05    3
 2.08548532e-08-4.68827401e-12-1.66736094e+04 2.02794895e+01                   4
CH3O2                   C   1H   3O   2     G    300.00   3500.00 1800.00      1
 5.64141817e+00 8.74328281e-03-3.21961406e-06 5.43695218e-10-3.45015008e-14    2
-1.19010148e+03-3.41914683e+00 1.44289632e+00 1.80733314e-02-1.09946545e-05    3
 3.42333984e-09-4.34452142e-13 3.21366390e+02 1.93041293e+01                   4
CH3OH                   C   1H   4O   1     G    300.00   3500.00 1800.00      1
 2.71701530e+00 1.21538353e-02-5.02107031e-06 1.01068070e-09-8.18460823e-14    2
-2.57693409e+04 9.47420540e+00 8.47330479e-01 1.63086904e-02-8.48344961e-06    3
 2.29304341e-09-2.59952013e-13-2.50962544e+04 1.95933297e+01                   4
CH3O                    C   1H   3O   1     G    300.00   3500.00 1740.00      1
 5.72238062e+00 5.90227637e-03-1.80340720e-06 2.13335009e-10-5.61816409e-15    2
-7.86252225e+01-7.49173677e+00 8.89660985e-01 1.70119767e-02-1.13807351e-05    3
 3.88280928e-09-5.32841479e-13 1.60316121e+03 1.85001134e+01                   4
CH2OH                   C   1H   3O   1     G    300.00   3500.00 1360.00      1
 5.04534950e+00 6.02727059e-03-2.11386821e-06 3.36085905e-10-2.00987482e-14    2
-4.03584143e+03-1.57524073e+00 2.34821579e+00 1.39600168e-02-1.08632206e-05    3
 4.62498416e-09-8.08499162e-13-3.30222106e+03 1.22661977e+01                   4
CH2O                    C   1H   2O   1     G    300.00   3500.00  700.00      1
 1.33335652e+00 1.00905183e-02-5.12952562e-06 1.25425207e-09-1.19639109e-13    2
-1.39080170e+04 1.59916144e+01 4.32621296e+00-7.01151853e-03 3.15176961e-05    3
-3.36478638e-08 1.23454023e-11-1.43270169e+04 2.62028902e+00                   4
HCO                     C   1H   1O   1     G    200.00   3500.00  770.00      1
 2.60049318e+00 5.29278258e-03-2.69184211e-06 7.21357798e-10-7.43521409e-14    2
 4.05725330e+03 1.07450933e+01 4.03483979e+00-2.15836864e-03 1.18233875e-05    3
-1.18459406e-08 4.00593954e-12 3.83636392e+03 4.20008770e+00                   4
HO2CHO                  C   1H   2O   3     G    300.00   3500.00 1750.00      1
 1.00230825e+01 4.43559488e-03-1.56185338e-06 2.43413972e-10-1.38379570e-14    2
-3.81313380e+04-2.33591553e+01 2.47434345e+00 2.16898555e-02-1.63512196e-05    3
 5.87745825e-09-8.18701426e-13-3.54892793e+04 1.72835404e+01                   4
HOCHO                   H   2C   1O   2     G    200.00   3500.00 1800.00      1
 3.79473661e+00 8.42765725e-03-3.84722250e-06 8.63389842e-10-7.73674422e-14    2
-4.73118221e+04 5.12933885e+00 1.85206266e+00 1.27447105e-02-7.44476686e-06    3
 2.19581368e-09-2.62426309e-13-4.66124595e+04 1.56434956e+01                   4
OCHO                    C   1O   2H   1     G    200.00   3500.00  700.00      1
 2.58373953e+00 8.99565940e-03-4.55939787e-06 1.11902584e-09-1.07899898e-13    2
-1.67164582e+04 1.34890938e+01 4.25809175e+00-5.72067562e-04 1.59428742e-05    3
-1.84069475e-08 6.86566202e-12-1.69508675e+04 6.00851172e+00                   4
C2H6                    C   2H   6          G    300.00   3500.00 1800.00      1
 4.07959141e+00 1.57445261e-02-5.96197393e-06 1.06867182e-09-7.61012340e-14    2
-1.25948053e+04-1.43089412e+00-2.41778724e-01 2.53475709e-02-1.39645112e-05    3
 4.03257452e-09-4.87754387e-13-1.10391121e+04 2.19572625e+01                   4
C2H5                    C   2H   5          G    300.00   3500.00 1800.00      1
 5.19791360e+00 1.11042800e-02-3.71281686e-06 5.47665571e-10-2.89412604e-14    2
 1.17176215e+04-4.91382513e+00 6.75421801e-01 2.11542617e-02-1.20878017e-05    3
 3.64951180e-09-4.59753237e-13 1.33457186e+04 1.95628439e+01                   4
C2H5O2H                 C   2H   6O   2     G    300.00   3500.00 1450.00      1
 1.00876750e+01 1.40221806e-02-4.79128015e-06 7.15474133e-10-3.78163629e-14    2
-2.40669299e+04-2.56733582e+01-5.77204918e-01 4.34425389e-02-3.52261336e-05    3
 1.47085102e-08-2.45040879e-12-2.09741147e+04 2.97412031e+01                   4
C2H5O2                  C   2H   5O   2     G    300.00   3500.00 1480.00      1
 9.29919683e+00 1.29334624e-02-4.54028592e-06 7.01327861e-10-3.92078228e-14    2
-7.64002445e+03-2.14311736e+01 2.00183268e-01 3.75253910e-02-2.94645378e-05    3
 1.19284684e-08-1.93568426e-12-4.94671644e+03 2.60335034e+01                   4
C2H4                    C   2H   4          G    300.00   3500.00 1650.00      1
 4.60402718e+00 9.50595350e-03-3.15129261e-06 4.53052074e-10-2.23949159e-14    2
 3.97229102e+03-3.77420905e+00-6.02932450e-02 2.08133970e-02-1.34307867e-05    3
 4.60638301e-09-6.51687481e-13 5.51151676e+03 2.10642172e+01                   4
C2H3                    C   2H   3          G    300.00   3500.00 1450.00      1
 4.18728376e+00 7.47581588e-03-2.58984227e-06 4.05265795e-10-2.35022721e-14    2
 3.38403785e+04 1.51958751e+00 1.23421214e+00 1.56222204e-02-1.10171572e-05    3
 4.27989337e-09-6.91541509e-13 3.46967692e+04 1.68637048e+01                   4
C2H2                    C   2H   2          G    300.00   3500.00  790.00      1
 4.37267454e+00 5.47212830e-03-2.03181542e-06 3.75019116e-10-2.77049062e-14    2
 2.58626597e+04-2.43835921e+00 7.70536907e-01 2.37107998e-02-3.66622044e-05    3
 2.95989761e-08-9.27579255e-12 2.64317975e+04 1.40907683e+01                   4
C2H                     C   2H   1          G    300.00   3500.00 1710.00      1
 3.41788257e+00 4.21328989e-03-1.58936946e-06 2.68739191e-10-1.73346359e-14    2
 6.72874491e+04 5.32512367e+00 4.60873599e+00 1.42766785e-03 8.54158643e-07    3
-6.83903344e-10 1.21940589e-13 6.68801772e+04-1.05894068e+00                   4
C2H5OH                  C   2H   6O   1     G    300.00   3500.00 1580.00      1
 7.32490827e+00 1.39762977e-02-4.67366748e-06 6.82063684e-10-3.47025038e-14    2
-3.18909574e+04-1.38313071e+01-4.22291411e-01 3.35894614e-02-2.32937596e-05    3
 8.53864266e-09-1.27783209e-12-2.94428423e+04 2.70882146e+01                   4
C2H5O                   C   2H   5O   1     G    300.00   3500.00  700.00      1
 1.68957255e+00 2.35453825e-02-1.23415273e-05 3.08911893e-09-2.98016648e-13    2
-3.10347953e+03 1.69410913e+01 3.27852943e+00 1.44656289e-02 7.11508755e-06    3
-1.54409905e-08 6.31987957e-12-3.32593350e+03 9.84203392e+00                   4
PC2H4OH                 C   2H   5O   1     G    300.00   3500.00 1470.00      1
 7.18479680e+00 1.17471700e-02-4.06239751e-06 6.31554725e-10-3.61645074e-14    2
-6.24418450e+03-9.60110092e+00 1.82077785e+00 2.63431399e-02-1.89562444e-05    3
 7.38613379e-09-1.18490244e-12-4.66716293e+03 1.83437446e+01                   4
SC2H4OH                 C   2H   5O   1     G    300.00   3500.00 1500.00      1
 6.63757422e+00 1.19924585e-02-4.07718738e-06 6.22004997e-10-3.47508084e-14    2
-9.66525354e+03-7.65007787e+00 1.23305393e+00 2.64045127e-02-1.84892415e-05    3
 7.02736239e-09-1.10231037e-12-8.04389745e+03 2.06149529e+01                   4
C2H4O2H                 C   2H   5O   2     G    300.00   3500.00 1440.00      1
 9.66417632e+00 1.29483231e-02-4.44318337e-06 6.83406482e-10-3.84804393e-14    2
 1.86599132e+03-2.38806241e+01 2.23212418e+00 3.35929124e-02-2.59479639e-05    3
 1.06393234e-08-1.76693824e-12 4.00642234e+03 1.46847781e+01                   4
C2H4O1-2                C   2H   4O   1     G    300.00   3500.00 1520.00      1
 6.04215804e+00 1.11433647e-02-3.80167462e-06 5.65226940e-10-2.94248186e-14    2
-9.44151524e+03-1.02352918e+01-2.19672856e+00 3.28246452e-02-2.51976751e-05    3
 9.94943769e-09-1.57288053e-12-6.93689371e+03 3.29622805e+01                   4
C2H3O1-2                C   2H   3O   1     G    200.00   3500.00 1800.00      1
 7.60993625e+00 6.11300596e-03-1.59366937e-06 1.28294159e-10 2.98968068e-15    2
 1.61313302e+04-1.70584528e+01 7.34197746e-02 2.28608204e-02-1.55501814e-05    3
 5.29737268e-09-7.14937891e-13 1.88444761e+04 2.37307466e+01                   4
CH3CHO                  C   2H   4O   1     G    300.00   3500.00 1800.00      1
 6.22195371e+00 1.06589270e-02-3.75190329e-06 6.00731628e-10-3.66603824e-14    2
-2.30621355e+04-8.31408577e+00 9.75916637e-01 2.23167871e-02-1.34667868e-05    3
 4.19883662e-09-5.36397187e-13-2.11735621e+04 2.00785613e+01                   4
CH3CO                   C   2H   3O   1     G    300.00   3500.00 1800.00      1
 6.07689016e+00 8.12979339e-03-2.81854999e-06 4.38698307e-10-2.55171837e-14    2
-4.06801047e+03-6.15492453e+00 1.47388064e+00 1.83587034e-02-1.13426417e-05    3
 3.59576931e-09-4.63999267e-13-2.41092705e+03 1.87575232e+01                   4
CH2CHO                  C   2H   3O   1     G    300.00   3500.00 1340.00      1
 6.47703792e+00 7.91358604e-03-2.83605891e-06 4.62112655e-10-2.83231297e-14    2
-1.16170812e+03-8.37157286e+00 7.37868281e-01 2.50454357e-02-2.20135026e-05    3
 1.00031294e-08-1.80836357e-12 3.76389339e+02 2.09962837e+01                   4
CH2CO                   C   2H   2O   1     G    300.00   3500.00 1360.00      1
 5.69523628e+00 6.46841658e-03-2.33588414e-06 3.83408110e-10-2.36897850e-14    2
-8.05944305e+03-4.61154403e+00 2.49503978e+00 1.58807592e-02-1.27171444e-05    3
 5.47226119e-09-9.59140718e-13-7.18898960e+03 1.18115657e+01                   4
HCCO                    C   2H   1O   1     G    300.00   3500.00 1220.00      1
 5.81420513e+00 3.89116779e-03-1.41168608e-06 2.35668533e-10-1.49424971e-14    2
 1.94026782e+04-4.94089647e+00 3.33028661e+00 1.20351629e-02-1.14247949e-05    3
 5.70731267e-09-1.13618105e-12 2.00087543e+04 7.53650387e+00                   4
HCOOH                   C   1H   2O   2     G    300.00   3500.00 1640.00      1
 5.21581644e+00 5.48253641e-03-1.72756111e-06 2.25438490e-10-8.81949912e-15    2
-4.56198641e+04-2.59494560e+00 1.19691275e+00 1.52847405e-02-1.06929917e-05    3
 3.86992247e-09-5.64381082e-13-4.43016637e+04 1.87820781e+01                   4
CH3CO3                  C   2H   3O   3     G    300.00   3500.00 1760.00      1
 1.40469381e+01 2.48483420e-03 1.65900439e-06-8.55133989e-10 9.82287244e-14    2
-2.73756816e+04-4.36816973e+01 2.64892548e+00 2.83894083e-02-2.04187576e-05    3
 7.50765465e-09-1.08966739e-12-2.33635811e+04 1.77505788e+01                   4
CH3CO3H                 C   2H   4O   3     G    300.00   3500.00 1240.00      1
 1.23807018e+01 1.08772145e-02-4.04888397e-06 6.94756696e-10-4.56573670e-14    2
-7.51809422e+04-3.74730276e+01-2.33886892e+00 5.83597007e-02-6.14873753e-05    3
 3.15756660e-08-6.27164715e-12-7.15304886e+04 3.67067395e+01                   4
CH2OHCHO                C   2H   4O   2     G    300.00   3500.00 1800.00      1
 8.91045186e+00 9.14305837e-03-2.53718677e-06 2.39203912e-10 8.50819938e-16    2
-4.09945450e+04-1.84179622e+01 1.56305396e+00 2.54706093e-02-1.61434792e-05    3
 5.27857147e-09-6.99061342e-13-3.83494818e+04 2.13476880e+01                   4
CHOCHO                  C   2H   2O   2     G    300.00   3500.00 1570.00      1
 9.97760259e+00 4.26981223e-03-1.12729433e-06 7.37809055e-11 5.98360578e-15    2
-2.96900177e+04-2.75230973e+01 7.08345765e-01 2.78857532e-02-2.36902952e-05    3
 9.65467301e-09-1.51963616e-12-2.67794711e+04 2.13768445e+01                   4
O2C2H4O2H               C   2H   5O   4     G    300.00   3500.00 1800.00      1
 1.24323243e+01 1.62358927e-02-6.84260319e-06 1.39267431e-09-1.12911127e-13    2
-1.87641105e+04-2.90906767e+01 5.81911522e+00 3.09319128e-02-1.90892866e-05    3
 5.92848299e-09-7.42884555e-13-1.63833552e+04 6.70139035e+00                   4
HO2CH2CHO               C   2H   4O   3     G    300.00   3500.00 1240.00      1
 1.23807018e+01 1.08772145e-02-4.04888397e-06 6.94756696e-10-4.56573670e-14    2
-7.51809422e+04-3.74730276e+01-2.33886892e+00 5.83597007e-02-6.14873753e-05    3
 3.15756660e-08-6.27164715e-12-7.15304886e+04 3.67067395e+01                   4
CH3OCHO                 C   2H   4O   2     G    300.00   3500.00  700.00      1
 5.02910657e+00-2.87377519e-02 6.15808970e-05-2.98073518e-08 4.29774802e-12    2
-4.07046731e+04 1.82412181e+01 2.12034974e-07-1.31715123e-09 2.87530013e-12    3
 2.88411189e-08-1.66481344e-11-4.00005982e+04 4.07099930e+01                   4
CH3OCO                  C   2H   3O   2     G    300.00   3500.00  730.00      1
 2.57527318e+00 2.11166692e-02-1.20149822e-05 3.14849390e-09-3.11411020e-13    2
-2.07588781e+04 1.60124236e+01 4.66126893e+00 9.68655552e-03 1.14715528e-05    3
-1.83003965e-08 7.03409940e-12-2.10634335e+04 6.60518516e+00                   4
C3H8                    C   3H   8          G    300.00   3500.00 1690.00      1
 8.33847007e+00 1.79340922e-02-5.80534981e-06 7.91037708e-10-3.43401227e-14    2
-1.70816233e+04-2.27461799e+01-1.38651266e+00 4.09518028e-02-2.62352705e-05    3
 8.85017800e-09-1.22652064e-12-1.37945792e+04 2.92742161e+01                   4
IC3H7                   C   3H   7          G    300.00   3500.00 1800.00      1
 6.05951251e+00 1.82035621e-02-6.54041321e-06 1.09272144e-09-7.13189353e-14    2
 7.29671818e+03-6.80793083e+00-6.08211221e-01 3.30207259e-02-1.88880497e-05    3
 5.66592015e-09-7.06485424e-13 9.69709872e+03 2.92791809e+01                   4
NC3H7                   C   3H   7          G    300.00   3500.00 1590.00      1
 7.21724982e+00 1.65877265e-02-5.58902439e-06 8.31338515e-10-4.40999325e-14    2
 8.50975633e+03-1.26938767e+01-1.37086178e-01 3.50892007e-02-2.30432453e-05    3
 8.14967015e-09-1.19478101e-12 1.08484352e+04 2.61969991e+01                   4
C3H6                    C   3H   6          G    298.00   3500.00 1800.00      1
 6.31755201e+00 1.65820017e-02-6.59972302e-06 1.29512916e-09-1.03784375e-13    2
-3.79456071e+02-1.05616187e+01-8.55987188e-02 3.08112255e-02-1.84574096e-05    3
 5.68686491e-09-7.13747674e-13 1.92567819e+03 2.40935687e+01                   4
CH2CHCH2                C   3H   5          G    298.00   3500.00 1600.00      1
 8.53877792e+00 1.04611885e-02-3.15379708e-06 3.85306884e-10-1.26413689e-14    2
 1.71766363e+04-2.28181758e+01-3.57888096e-01 3.27028536e-02-2.40053580e-05    3
 9.07345729e-09-1.37016487e-12 2.00235695e+04 2.42845603e+01                   4
C3H5-S                  C   3H   5          G    300.00   3500.00 1800.00      1
 6.52599516e+00 1.37686655e-02-5.50691342e-06 1.07278366e-09-8.39560017e-14    2
 2.86430050e+04-9.99635700e+00 1.54227621e+00 2.48435965e-02-1.47360226e-05    3
 4.49097224e-09-5.58704416e-13 3.04371438e+04 1.69765696e+01                   4
C3H5-T                  C   3H   5          G    300.00   3500.00  770.00      1
 1.49331935e+00 2.33788729e-02-1.18550710e-05 2.86552470e-09-2.68203790e-13    2
 2.87117775e+04 1.76892214e+01 2.52238869e+00 1.80330581e-02-1.44114618e-06    3
-6.15086046e-09 2.65919399e-12 2.85533009e+04 1.29935191e+01                   4
C3H5O                   C   3H   5O   1     G    300.00   3500.00 1610.00      1
 9.11079978e+00 1.37589661e-02-5.15319199e-06 9.32421983e-10-6.74695911e-14    2
 7.77376170e+03-2.10036658e+01 9.27196847e-01 3.40908988e-02-2.40959865e-05    3
 8.77622923e-09-1.28545208e-12 1.04088818e+04 2.23747992e+01                   4
C3H6O                   C   3H   6O   1     G    300.00   3500.00 1550.00      1
 9.00938222e+00 1.57632590e-02-5.29374355e-06 7.64253417e-10-3.74126438e-14    2
-1.56669515e+04-2.44960178e+01-1.88321638e+00 4.38731909e-02-3.24969034e-05    3
 1.24645372e-08-1.92455519e-12-1.22902459e+04 3.28282089e+01                   4
CH3CHCHO                C   3H   5O   1     G    300.00   3500.00 1800.00      1
 6.70347362e+00 1.89922318e-02-9.18109977e-06 2.14445657e-09-1.96154637e-13    2
-6.21094363e+03-1.05801331e+01 2.92067498e-01 3.32398010e-02-2.10540741e-05    3
 6.54185446e-09-8.06904344e-13-3.90283743e+03 2.41197343e+01                   4
AC4H7OOH                C   4H   8O   2     G    300.00   3500.00 1660.00      1
 1.22738272e+01 2.55483383e-02-9.81265077e-06 1.82078670e-09-1.35039880e-13    2
-1.24525960e+04-3.36837474e+01 1.60151447e+00 5.12647544e-02-3.30503762e-05    3
 1.11532065e-08-1.54052480e-12-8.90938817e+03 2.32129081e+01                   4
CH3CHCO                 C   3H   4O   1     G    300.00   3500.00 1280.00      1
 6.99681463e+00 1.49445085e-02-6.71568578e-06 1.45955079e-09-1.25293200e-13    2
-1.29366480e+04-1.07908059e+01 1.50068777e+00 3.21199049e-02-2.68431035e-05    3
 1.19425808e-08-2.17276001e-12-1.15296395e+04 1.70816035e+01                   4
AC3H5OOH                C   3H   6O   2     G    298.00   3500.00 1800.00      1
 1.36957657e+01 1.27112963e-02-4.21186263e-06 6.49030109e-10-3.94931202e-14    2
-1.11479407e+04-4.31791016e+01 4.22354618e+00 3.37606729e-02-2.17530098e-05    3
 7.14575129e-09-9.41815506e-13-7.73794171e+03 8.08652616e+00                   4
C3H6OH1-2               C   3H   7O   1     G    300.00   3500.00 1800.00      1
 8.46016352e+00 1.89669003e-02-7.38013554e-06 1.39189577e-09-1.05413394e-13    2
-1.21581707e+04-1.51603324e+01 4.08605477e-01 3.68592515e-02-2.22904282e-05    3
 6.91422639e-09-8.72403758e-13-9.25960980e+03 2.84163793e+01                   4
C3H6OH2-1               C   3H   7O   1     G    300.00   3500.00 1590.00      1
 8.99548234e+00 1.75103792e-02-6.94615357e-06 1.37004323e-09-1.07539337e-13    2
-1.65436320e+04-1.93287236e+01 1.31207693e+00 3.68397010e-02-2.51813628e-05    3
 9.01583327e-09-1.30970758e-12-1.41003090e+04 2.13023225e+01                   4
HOC3H6O2                C   3H   7O   3     G    300.00   3500.00 1480.00      1
 1.24409055e+01 2.15172909e-02-8.97737594e-06 1.82414691e-09-1.48047122e-13    2
-3.10315628e+04-3.23089026e+01 2.93449048e+00 4.72103044e-02-3.50175923e-05    3
 1.35539741e-08-2.12943685e-12-2.82176640e+04 1.72809693e+01                   4
SC3H5OH                 C   3H   6O   1     G    300.00   3500.00 1260.00      1
 7.83167544e+00 1.85990426e-02-7.98421836e-06 1.67672190e-09-1.40411942e-13    2
-2.22362405e+04-1.56369776e+01-5.71229678e-02 4.36428470e-02-3.77982713e-05    3
 1.74513531e-08-3.27029908e-12-2.02482633e+04 2.42451084e+01                   4
C3H5OH                  C   3H   6O   1     G    300.00   3500.00 1630.00      1
 9.39463114e+00 1.51343106e-02-4.86246276e-06 6.64177249e-10-2.94552530e-14    2
-2.20582199e+04-2.45922026e+01 4.73537667e-01 3.70265645e-02-2.50087087e-05    3
 8.90395064e-09-1.29322418e-12-1.91499434e+04 2.28055845e+01                   4
CH2CCH2OH               C   3H   5O   1     G    300.00   3500.00 1800.00      1
 7.15397365e+00 1.62590933e-02-7.06959971e-06 1.52062107e-09-1.30983749e-13    2
 1.01359982e+04-8.36739478e+00 2.39300609e+00 2.68390212e-02-1.58862063e-05    3
 4.78603091e-09-5.84512894e-13 1.18499465e+04 1.73999548e+01                   4
PC3H4                   C   3H   4          G    300.00   3500.00 1570.00      1
 6.45797858e+00 1.06371316e-02-3.61161722e-06 5.39412691e-10-2.85851275e-14    2
 1.94136786e+04-1.10770989e+01 1.72714322e+00 2.26902153e-02-1.51273023e-05    3
 5.42930020e-09-8.07229635e-13 2.08991609e+04 1.38804115e+01                   4
AC3H4                   C   3H   4          G    300.00   3500.00 1420.00      1
 6.37608366e+00 1.10282079e-02-3.89476312e-06 6.16686076e-10-3.59564768e-14    2
 2.00917847e+04-1.13283006e+01 5.08248696e-01 2.75573205e-02-2.13550933e-05    3
 8.81402419e-09-1.47914981e-12 2.17582498e+04 1.90382079e+01                   4
C3H3                    C   3H   3          G    300.00   3500.00  840.00      1
 5.75057762e+00 1.05635747e-02-4.84060952e-06 1.09040068e-09-9.80036130e-14    2
 4.00565408e+04-5.04125059e+00 1.75584147e+00 2.95861278e-02-3.88094543e-05    3
 2.80498013e-08-8.12163476e-12 4.07276565e+04 1.35345464e+01                   4
C3H2                    C   3H   2          G    300.00   3500.00 1260.00      1
 6.42043189e+00 6.05128866e-03-2.30888141e-06 4.10631875e-10-2.84293474e-14    2
 6.08598164e+04-8.32404334e+00 2.15397882e+00 1.95955841e-02-1.84330427e-05    3
 8.94193413e-09-1.72114805e-12 6.19349626e+04 1.32451538e+01                   4
C2H5CHO                 C   3H   6O   1     G    300.00   3500.00 1710.00      1
 9.33264604e+00 1.46861072e-02-4.56011955e-06 5.69518135e-10-1.90908109e-14    2
-2.69164882e+04-2.52385565e+01-9.86882752e-02 3.67477080e-02-2.39124009e-05    3
 8.11426720e-09-1.12212430e-12-2.36909719e+04 2.53220280e+01                   4
CH2CH2CHO               C   3H   5O   1     G    300.00   3500.00  700.00      1
 1.38640400e+00 2.84363938e-02-1.56688640e-05 4.07196321e-09-4.03232083e-13    2
 6.14151634e+02 2.19844218e+01 2.41071832e+00 2.25831692e-02-3.12623980e-06    3
-7.87339320e-09 3.86296664e-12 4.70747631e+02 1.74080446e+01                   4
RALD3                   C   3H   5O   1     G    300.00   3500.00 1140.00      1
-6.08013768e+00 4.60180078e-02-2.61696720e-05 6.65382129e-09-6.35305357e-13    2
-2.14966001e+03 5.90959840e+01 7.04072886e+00-2.01204450e-05 3.44068124e-05    3
-2.87710234e-08 7.13330094e-12-5.14121758e+03-5.92381685e+00                   4
C2H3CHO                 C   3H   4O   1     G    300.00   3500.00 1600.00      1
 9.22597839e+00 1.12038372e-02-3.67974365e-06 5.08180252e-10-2.25803375e-14    2
-1.23719484e+04-2.08137560e+01 8.18908043e-01 3.22215131e-02-2.33838148e-05    3
 8.71820989e-09-1.30539747e-12-9.68168587e+03 2.36968522e+01                   4
CH3COCH3                C   3H   6O   1     G    300.00   3500.00 1790.00      1
 9.79507855e+00 1.35932465e-02-4.01642284e-06 4.43034305e-10-7.94380246e-15    2
-3.07542949e+04-2.70699391e+01-7.54581368e-03 3.54985524e-02-2.23728244e-05    3
 7.27968292e-09-9.62782995e-13-2.72449554e+04 2.59292980e+01                   4
CH3COCH2                C   3H   5O   1     G    300.00   3500.00 1590.00      1
 8.40473847e+00 1.29432044e-02-4.25667366e-06 6.02254911e-10-2.86748418e-14    2
-7.89528923e+03-1.63899805e+01 1.00367440e+00 3.15622335e-02-2.18217955e-05    3
 7.96708586e-09-1.18666713e-12-5.54175085e+03 2.27480006e+01                   4
NC4H10                  C   4H  10          G    300.00   3500.00 1800.00      1
 1.54355362e+01 1.56272553e-02-3.14851999e-06-5.94424210e-11 5.32964638e-14    2
-2.28455262e+04-6.02417835e+01-1.20836758e+00 5.26137081e-02-3.39705640e-05    3
 1.13561294e-08-1.53219963e-12-1.68537208e+04 2.98384958e+01                   4
PC4H9                   C   4H   9          G    300.00   3500.00  950.00      1
 3.94763006e+00 3.16286394e-02-1.12984867e-05 1.11637450e-09 5.54031605e-14    2
 6.05554723e+03 7.76350061e+00-2.76188385e-01 4.94131381e-02-3.93792741e-05    3
 2.08221903e-08-5.13033783e-12 6.85807273e+03 2.79243295e+01                   4
SC4H9                   C   4H   9          G    300.00   3500.00  850.00      1
 3.40122928e+00 3.20901863e-02-1.12255470e-05 9.71712110e-10 8.30726274e-14    2
 4.66283101e+03 1.05291639e+01 2.36336421e-01 4.69837998e-02-3.75083943e-05    3
 2.15857099e-08-5.97986791e-12 5.20086280e+03 2.52835874e+01                   4
IC4H10                  C   4H  10          G    300.00   3500.00 1260.00      1
 5.51955795e+00 3.23747266e-02-1.18655436e-05 1.37455177e-09 1.57073481e-14    2
-1.97025810e+04-6.34483426e+00-1.85965329e+00 5.58007941e-02-3.97537191e-05    3
 1.61302002e-08-2.91200067e-12-1.78430198e+04 3.09610166e+01                   4
IC4H9                   C   4H   9          G    300.00   3500.00 1430.00      1
 7.95880517e+00 2.55088283e-02-8.62221490e-06 8.09648920e-10 4.02033223e-14    2
 3.37759297e+03-1.61084037e+01-1.15582377e+00 5.10042938e-02-3.53657102e-05    3
 1.32774789e-08-2.13948724e-12 5.98437685e+03 3.11244820e+01                   4
TC4H9                   C   4H   9          G    300.00   3500.00 1400.00      1
 7.90871689e+00 2.55264450e-02-8.65284049e-06 8.24419700e-10 3.80550657e-14    2
 8.35470579e+02-1.73299272e+01-1.29900233e+00 5.18342142e-02-3.68397361e-05    3
 1.42467509e-08-2.35878980e-12 3.41363196e+03 3.01901373e+01                   4
IC4H8                   C   4H   8          G    300.00   3500.00 1800.00      1
 7.63433967e+00 2.47722696e-02-1.05415828e-05 2.18152373e-09-1.80119594e-13    2
-6.21385767e+03-1.72949366e+01 7.17301599e-01 4.01434653e-02-2.33509125e-05    3
 6.92571993e-09-8.39035733e-13-3.72372397e+03 2.01415164e+01                   4
IC4H7                   C   4H   7          G    300.00   3500.00  700.00      1
 1.18177117e+00 3.67769037e-02-1.77031337e-05 3.74786266e-09-2.92191284e-13    2
 1.31214242e+04 2.00120540e+01 3.86130010e+00 2.14653098e-02 1.51074247e-05    3
-2.75002882e-08 1.08678626e-11 1.27462902e+04 8.04059663e+00                   4
IC4H7O                  C   4H   7O   1     G    300.00   3500.00 1800.00      1
 1.18822163e+01 1.89918532e-02-7.42296498e-06 1.41442848e-09-1.08683660e-13    2
 1.15971319e+03-3.56333819e+01 1.50010972e+00 4.20632012e-02-2.66490883e-05    3
 8.53521488e-09-1.09768177e-12 4.89727156e+03 2.05567447e+01                   4
C4H8-1                  C   4H   8          G    300.00   3500.00 1800.00      1
 1.03330449e+01 1.99470428e-02-7.40538998e-06 1.30472507e-09-9.09598189e-14    2
-5.56551437e+03-3.07722296e+01-6.91489888e-01 4.44460090e-02-2.78211951e-05    3
 8.86613439e-09-1.14115556e-12-1.59668184e+03 2.88948525e+01                   4
C4H8-2                  C   4H   8          G    300.00   3500.00 1800.00      1
 5.15907399e+00 2.89997694e-02-1.32974598e-05 2.96139017e-09-2.60424474e-13    2
-4.76704683e+03-3.39008062e+00 5.60608454e-01 3.92185817e-02-2.18131368e-05    3
 6.11534459e-09-6.98473698e-13-3.11159924e+03 2.14977742e+01                   4
C4H71-3                 C   4H   7          G    300.00   3500.00 1420.00      1
 8.33017754e+00 1.98466503e-02-6.37614061e-06 5.28652768e-10 3.81103734e-14    2
 1.19533850e+04-1.83767119e+01-1.12550124e+00 4.64823652e-02-3.45124591e-05    3
 1.37381920e-08-2.28751273e-12 1.46387978e+04 3.05571711e+01                   4
C4H71-4                 C   4H   7          G    300.00   3500.00 1530.00      1
 8.45916998e+00 1.93968541e-02-5.99075605e-06 3.82147970e-10 5.73994809e-14    2
 1.98988324e+04-1.80212793e+01-3.29329052e-01 4.23733221e-02-2.85167051e-05    3
 1.01973763e-08-1.54639600e-12 2.25881131e+04 2.81156134e+01                   4
C4H71-O                 C   4H   7O   1     G    300.00   3500.00 1600.00      1
 1.37371777e+01 1.70982846e-02-6.55972544e-06 1.21466090e-09-8.98269615e-14    2
-3.28789072e+01-4.64105970e+01-1.48200925e+00 5.51462520e-02-4.22296948e-05    3
 1.60771481e-08-2.41209059e-12 4.83726091e+03 3.41662556e+01                   4
C4H6                    C   4H   6          G    200.00   3500.00 1800.00      1
 9.30872521e+00 1.50139591e-02-5.06688177e-06 7.84148097e-10-4.70262839e-14    2
 8.60829987e+03-2.47389586e+01 4.65225109e-01 3.46661815e-02-2.14437338e-05    3
 6.84964885e-09-8.89456944e-13 1.17919599e+04 2.31239087e+01                   4
C4H5                    C   4H   5          G    300.00   3500.00 1800.00      1
 1.90192654e+01-1.91794386e-03 4.88814514e-06-1.91833948e-09 2.24139237e-13    2
 3.48592740e+04-7.70423351e+01-2.01742308e-01 4.07954066e-02-3.07063136e-05    3
 1.12647934e-08-1.60685144e-12 4.17788367e+04 2.69857683e+01                   4
C4H4                    C   4H   4          G    300.00   3500.00 1290.00      1
 7.65777119e+00 1.26498258e-02-4.62248950e-06 7.81217082e-10-5.07629107e-14    2
 3.13366016e+04-1.49692661e+01 7.13119716e-01 3.41836288e-02-2.96617954e-05    3
 1.37214268e-08-2.55855550e-12 3.31283217e+04 2.03030643e+01                   4
C4H3                    C   4H   3          G    300.00   3500.00 1590.00      1
 1.30208969e+01 1.53590364e-03 1.80568200e-06-9.30237204e-10 1.18077198e-13    2
 6.01811751e+04-4.25791500e+01 2.34662666e+00 2.83894138e-02-2.35278181e-05    3
 9.69177543e-09-1.55205057e-12 6.35755930e+04 1.38680560e+01                   4
C4H2                    C   4H   2          G    300.00   3500.00  720.00      1
 7.13414735e+00 1.00526308e-02-4.84819206e-06 1.14884604e-09-1.07722834e-13    2
 5.27577824e+04-1.36443516e+01-4.34754087e-01 5.21020832e-02-9.24512179e-05    3
 8.22627589e-08-2.82722759e-11 5.38477042e+04 2.03848077e+01                   4
C6H6                    C   6H   6          G    300.00   3500.00 1410.00      1
 1.15055544e+01 1.99961045e-02-7.07935460e-06 1.10673028e-09-6.24178899e-14    2
 4.11452290e+03-4.24445091e+01-6.99882110e+00 7.24907868e-02-6.29247613e-05    3
 2.75111779e-08-4.74405754e-12 9.33275680e+03 5.31863191e+01                   4
FULVENE                 C   6H   6          G    200.00   3500.00 1560.00      1
 1.44152220e+01 1.47750067e-02-3.90939181e-06 2.82308156e-10 1.62511622e-14    2
 1.91167581e+04-5.54965184e+01-3.67012639e+00 6.11476948e-02-4.84985149e-05    3
 1.93374890e-08-3.03746371e-12 2.47593868e+04 3.97971310e+01                   4
C6H5                    C   6H   5          G    300.00   3500.00 1390.00      1
 1.12331261e+01 1.77269649e-02-6.33615682e-06 1.00236865e-09-5.75481750e-14    2
 3.49856300e+04-3.80075865e+01-6.76261385e+00 6.95132669e-02-6.22206553e-05    3
 2.78054854e-08-4.87825263e-12 3.99884457e+04 5.47375207e+01                   4
C5H6                    C   5H   6          G    200.00   3500.00 1630.00      1
 1.35786764e+01 1.28174257e-02-3.11961936e-06 1.29368393e-10 2.76958521e-14    2
 9.43770579e+03-5.26289052e+01-4.05866643e+00 5.60992486e-02-4.29495178e-05    3
 1.64197154e-08-2.47082363e-12 1.51874796e+04 4.10783319e+01                   4
C5H5                    C   5H   5          G    300.00   3500.00  700.00      1
 4.01652588e+00 2.68451887e-02-1.26423015e-05 2.78092323e-09-2.35299425e-13    2
 2.91110159e+04 1.44025731e+00-2.58737467e+00 6.45817633e-02-9.35063898e-05    3
 7.97943407e-08-2.77400914e-11 3.00355619e+04 3.09448142e+01                   4
MCPTD                   C   6H   8          G    300.00   3500.00 1470.00      1
 1.21408016e+01 2.34281374e-02-7.98702759e-06 1.18908391e-09-6.20202054e-14    2
 7.23040214e+03-4.21606537e+01-5.49894699e+00 7.14274534e-02-5.69659215e-05    3
 2.34017342e-08-3.83968182e-12 1.24164882e+04 4.97368686e+01                   4
C10H8                   C  10H   8          G    300.00   3500.00 1370.00      1
 1.51184828e+01 3.89675576e-02-1.78248658e-05 3.92092279e-09-3.39215689e-13    2
 1.01121562e+04-6.09041102e+01-8.71832426e+00 1.08564074e-01-9.40254318e-05    3
 4.10014902e-08-7.10574258e-12 1.66434413e+04 6.15987877e+01                   4
NC3H7O2                 C   3H   7O   2     G    300.00   3500.00 1650.00      1
 9.25591855e+00 2.27563801e-02-9.54934453e-06 1.92559465e-09-1.53946670e-13    2
-9.34005086e+03-1.86388081e+01 1.92964396e+00 4.05170458e-02-2.56954042e-05    3
 8.44925513e-09-1.14238008e-12-6.92238025e+03 2.03750491e+01                   4
IC3H7O2                 C   3H   7O   2     G    300.00   3500.00 1260.00      1
 7.34738699e+00 2.68252330e-02-1.24179691e-05 2.76645854e-09-2.42147350e-13    2
-1.06484855e+04-8.92587195e+00 1.07341266e+00 4.67426118e-02-3.61291344e-05    3
 1.53120486e-08-2.73135173e-12-9.06744395e+03 2.27924165e+01                   4
C3H7OOH                 C   3H   8O   2     G    300.00   3500.00 1530.00      1
 1.13871492e+01 1.97925480e-02-6.62893779e-06 9.67106876e-10-4.94700798e-14    2
-2.73563036e+04-2.91104777e+01-9.73590405e-01 5.21082072e-02-3.83109566e-05    3
 1.47719081e-08-2.30515656e-12-2.35739173e+04 3.57795697e+01                   4
C3-OQOOH                C   3H   6O   3     G    300.00   3500.00 1350.00      1
 1.12132537e+01 2.34709018e-02-1.13098317e-05 2.59008079e-09-2.30885269e-13    2
-3.91289882e+04-2.66260028e+01 8.46220450e-01 5.41880374e-02-4.54399823e-05    3
 1.94444762e-08-3.35206960e-12-3.63298893e+04 2.65001343e+01                   4
CHOCH2CHO               C   3H   4O   2     G    300.00   3500.00 1370.00      1
 1.06304440e+01 1.18394227e-02-4.21486308e-06 6.67473434e-10-3.88516159e-14    2
-4.37970340e+04-2.83088260e+01-8.46550190e-01 4.53488948e-02-4.09040660e-05    3
 1.85211002e-08-3.29681270e-12-4.06523375e+04 3.06741176e+01                   4
CH2OHCH2CHO             C   3H   6O   2     G    300.00   3500.00 1800.00      1
 1.08721654e+01 1.63593216e-02-6.08637842e-06 1.10130849e-09-8.02911325e-14    2
-4.55272952e+04-2.70748520e+01 2.66105929e+00 3.46062241e-02-2.12921305e-05    3
 6.73306853e-09-8.62480026e-13-4.25712970e+04 1.73653673e+01                   4
CH3CO2H                 C   2H   4O   2     G    300.00   3500.00 1800.00      1
 1.06195365e+01 8.83226600e-03-2.54924379e-06 2.13473353e-10 7.27652554e-15    2
-5.71972759e+04-3.23726793e+01-7.52613551e-01 3.41037106e-02-2.36087809e-05    3
 8.01330193e-09-1.07603300e-12-5.31033019e+04 2.91757692e+01                   4
HCO3                    C   1H   1O   3     G    300.00   3500.00 1490.00      1
 7.67843584e+00 4.62692543e-03-1.54275270e-06 2.12409842e-10-8.98166116e-15    2
-1.61147276e+04-1.27152259e+01 2.31459990e+00 1.90264850e-02-1.60389536e-05    3
 6.69840577e-09-1.09723601e-12-1.45163044e+04 1.53011516e+01                   4
HCO3H                   C   1H   2O   3     G    300.00   3500.00 1750.00      1
 1.00230668e+01 4.43563253e-03-1.56188514e-06 2.43424395e-10-1.38391380e-14    2
-3.81313332e+04-2.33590722e+01 2.47434199e+00 2.16898607e-02-1.63512235e-05    3
 5.87745807e-09-8.18701091e-13-3.54892796e+04 1.72835470e+01                   4
CH2OHCOCH3              C   3H   6O   2     G    300.00   3500.00 1460.00      1
 1.16062110e+01 1.59761333e-02-5.42430575e-06 8.11522092e-10-4.31363774e-14    2
-4.81919050e+04-3.20429615e+01 9.15361352e-01 4.52661324e-02-3.55167705e-05    3
 1.45523736e-08-2.39602191e-12-4.50701769e+04 2.35800153e+01                   4
NC3-QOOH                C   3H   7O   2     G    300.00   3500.00 1800.00      1
 1.29748618e+01 1.76433870e-02-7.16935406e-06 1.42696153e-09-1.14477043e-13    2
-5.86411825e+03-3.67690498e+01 1.55643299e+00 4.30176732e-02-2.83145926e-05    3
 9.25853134e-09-1.20219507e-12-1.75348388e+03 2.50298688e+01                   4
IC3-QOOH                C   3H   7O   2     G    300.00   3500.00 1270.00      1
 1.04498043e+01 2.29490980e-02-1.05757759e-05 2.34172678e-09-2.03669154e-13    2
-5.22299426e+03-2.40008692e+01-1.71110877e-01 5.64007993e-02-5.00856593e-05    3
 2.30818230e-08-4.28636527e-12-2.52528181e+03 2.97774852e+01                   4
NC3-OOQOOH              C   3H   7O   4     G    300.00   3500.00 1260.00      1
 1.11683562e+01 2.95822139e-02-1.42526305e-05 3.27126849e-09-2.92476812e-13    2
-2.00281219e+04-2.06289848e+01 2.57588692e+00 5.68598942e-02-4.67260594e-05    3
 2.04529769e-08-3.70154594e-12-1.78628196e+04 2.28105329e+01                   4
IC3-OOQOOH              C   3H   7O   4     G    300.00   3500.00 1220.00      1
 1.23035624e+01 2.79964884e-02-1.33482910e-05 3.03524084e-09-2.69271163e-13    2
-2.25784829e+04-2.78550798e+01 1.73143844e+00 6.26591899e-02-5.59663668e-05    3
 2.63238068e-08-5.04151829e-12-1.99988847e+04 2.52515831e+01                   4
CH2COOH                 C   2H   3O   2     G    300.00   3500.00 1440.00      1
 1.01170850e+01 5.56298782e-03-8.24128628e-07-2.50442742e-11 1.25384218e-14    2
-3.40138321e+04-2.77197730e+01 4.26277933e-01 3.24818963e-02-2.88646583e-05    3
 1.29566824e-08-2.24123357e-12-3.12228797e+04 2.25664553e+01                   4
IC4-OQOOH               C   4H   8O   3     G    300.00   3500.00 1570.00      1
 1.51567879e+01 2.57227734e-02-1.11020451e-05 2.28943518e-09-1.86269530e-13    2
-4.30658407e+04-4.59845002e+01 9.69279338e-01 6.18692920e-02-4.56369355e-05    3
 1.69539322e-08-2.52138051e-12-3.86109630e+04 2.88616666e+01                   4
NC4-OQOOH               C   4H   8O   3     G    300.00   3500.00 1330.00      1
 1.18153445e+01 3.20093755e-02-1.53334982e-05 3.50316407e-09-3.12136547e-13    2
-4.27660549e+04-2.73083214e+01 2.51946601e+00 5.99669047e-02-4.68645461e-05    3
 1.93082006e-08-3.28300808e-12-4.02933512e+04 2.01899074e+01                   4
C4H9OOH                 C   4H  10O   2     G    300.00   3500.00 1780.00      1
 1.73966948e+01 2.30088698e-02-8.34646932e-06 1.39883190e-09-9.01677554e-14    2
-3.38614042e+04-6.23628946e+01 1.12895120e+00 5.95655969e-02-3.91527000e-05    3
 1.29367460e-08-1.71066131e-12-2.80700874e+04 2.54997628e+01                   4
C5EN-OQOOH-35           C   5H   8O   3     G    300.00   3500.00 1580.00      1
 1.69833146e+01 2.73095032e-02-1.19226853e-05 2.48166925e-09-2.03420392e-13    2
-3.51234520e+04-5.58041780e+01 1.44561329e+00 6.66454559e-02-4.92669442e-05    3
 1.82387405e-08-2.69662788e-12-3.02135384e+04 2.62635800e+01                   4
NC5H10-O                C   5H  10O   1     G    300.00   3500.00 1800.00      1
 1.40073101e+01 3.04405284e-02-1.35854526e-05 2.90305354e-09-2.44985844e-13    2
-2.55455866e+04-5.25239383e+01-3.79263098e+00 6.99959530e-02-4.65483064e-05    3
 1.51115179e-08-1.94060590e-12-1.91376078e+04 4.38130562e+01                   4
NC5-OQOOH               C   5H  10O   3     G    300.00   3500.00 1410.00      1
 1.42172630e+01 3.77707683e-02-1.76257936e-05 3.93443034e-09-3.43954252e-13    2
-4.65061050e+04-3.85369191e+01 2.52749929e+00 7.09332187e-02-5.29049961e-05    3
 2.06149043e-08-3.30148510e-12-4.32095916e+04 2.18759162e+01                   4
NC5H11OOH               C   5H  12O   2     G    300.00   3500.00 1630.00      1
 1.66988185e+01 3.44172712e-02-1.43139761e-05 2.85300849e-09-2.25350876e-13    2
-3.73755763e+04-5.75775302e+01 6.24289379e-02 7.52427671e-02-5.18834508e-05    3
 1.82188468e-08-2.58207455e-12-3.19521133e+04 3.08116402e+01                   4
NC4-QOOH                C   4H   9O   2     G    300.00   3500.00 1760.00      1
 1.83774568e+01 1.83354725e-02-6.23923380e-06 9.66797423e-10-5.61281944e-14    2
-1.29135491e+04-6.55986639e+01 1.19976578e+00 5.73756794e-02-3.95121374e-05    3
 1.35701700e-08-1.84637998e-12-6.86700189e+03 2.69845517e+01                   4
NC4H9-OO                C   4H   9O   2     G    300.00   3500.00 1320.00      1
 8.96630114e+00 3.41074657e-02-1.57641000e-05 3.50715782e-09-3.06662916e-13    2
-1.40847395e+04-1.58347447e+01 9.44281656e-01 5.84166156e-02-4.33881341e-05    3
 1.74586902e-08-2.94899859e-12-1.19669263e+04 2.50940293e+01                   4
IC4H9T-OO               C   4H   9O   2     G    300.00   3500.00 1260.00      1
 9.11667611e+00 3.41757258e-02-1.58797345e-05 3.54686464e-09-3.10976548e-13    2
-1.64591648e+04-1.96564028e+01 4.84069010e-01 6.15808277e-02-4.85048558e-05    3
 2.08088336e-08-3.73597039e-12-1.42837478e+04 2.39860330e+01                   4
IC4T-QOOH               C   4H   9O   2     G    300.00   3500.00 1270.00      1
 1.20890742e+01 3.03954175e-02-1.40883982e-05 3.13822121e-09-2.74437748e-13    2
-1.09705556e+04-3.28537329e+01-4.26302142e-01 6.98139255e-02-6.06456912e-05    3
 2.75777451e-08-5.08536764e-12-7.79165002e+03 3.05171096e+01                   4
IC4P-QOOH               C   4H   9O   2     G    300.00   3500.00 1350.00      1
 1.14809469e+01 3.08095616e-02-1.41939360e-05 3.14755455e-09-2.74422165e-13    2
-7.45268236e+03-2.80879239e+01-1.93281563e-01 6.53998681e-02-5.26276099e-05    3
 2.21271466e-08-3.78916143e-12-4.30064068e+03 3.17369695e+01                   4
IC4H9P-OO               C   4H   9O   2     G    300.00   3500.00 1380.00      1
 8.54295826e+00 3.45220773e-02-1.59311943e-05 3.53852672e-09-3.08950056e-13    2
-1.29532173e+04-1.39825068e+01 7.00555203e-01 5.72536803e-02-4.06394585e-05    3
 1.54748862e-08-2.47133403e-12-1.07887140e+04 2.63784632e+01                   4
NC4-OOQOOH              C   4H   9O   4     G    300.00   3500.00 1230.00      1
 1.51474113e+01 3.37812811e-02-1.58996825e-05 3.57608795e-09-3.14486518e-13    2
-2.85698876e+04-4.24732202e+01 1.10123476e+00 7.94599040e-02-7.16053202e-05    3
 3.37688455e-08-6.45122585e-12-2.51145282e+04 2.81992196e+01                   4
IC4T-OOQOOH             C   4H   9O   4     G    300.00   3500.00 1240.00      1
 1.39939782e+01 3.54845223e-02-1.68915059e-05 3.83671077e-09-3.40131615e-13    2
-2.83614519e+04-3.70531088e+01 1.55094394e+00 7.56233423e-02-6.54465302e-05    3
 2.99415625e-08-5.60320657e-12-2.52755794e+04 2.56539769e+01                   4
IC4P-OOQOOH             C   4H   9O   4     G    300.00   3500.00 1290.00      1
 1.30518446e+01 3.65484801e-02-1.74274782e-05 3.96741951e-09-3.52552034e-13    2
-2.47096139e+04-3.04334702e+01 1.64511787e+00 7.19181753e-02-5.85550308e-05    3
 2.52219687e-08-4.47165071e-12-2.17666784e+04 2.75020267e+01                   4
C5EN-QOOH               C   5H   9O   2     G    300.00   3500.00 1420.00      1
 1.28791275e+01 3.32930454e-02-1.55378924e-05 3.46674396e-09-3.02869803e-13    2
 3.23011716e+03-3.38507184e+01 1.34404411e+00 6.57862381e-02-4.98616876e-05    3
 1.95812018e-08-3.13992224e-12 6.50608085e+03 2.58442475e+01                   4
C5EN-OO                 C   5H   9O   2     G    300.00   3500.00 1280.00      1
 1.00840321e+01 3.69913036e-02-1.74216180e-05 3.93130749e-09-3.47257402e-13    2
-8.98415155e+02-1.96513637e+01 4.09897282e-01 6.72229749e-02-5.28493577e-05    3
 2.23832553e-08-3.95115346e-12 1.57816336e+03 2.94089022e+01                   4
C5EN-OOQOOH-35          C   5H   9O   4     G    300.00   3500.00 1160.00      1
 1.36699765e+01 4.21231934e-02-2.15503712e-05 5.21806335e-09-4.87293013e-13    2
-1.42354804e+04-3.35883365e+01 5.24578569e-01 8.74521518e-02-8.01654036e-05    3
 3.89048636e-08-7.74737927e-12-1.11857480e+04 3.17816498e+01                   4
NC5H12OO                C   5H  11O   2     G    300.00   3500.00 1300.00      1
 1.06544848e+01 4.16170555e-02-1.93382868e-05 4.32113942e-09-3.79088223e-13    2
-1.98652039e+04-2.50234586e+01 3.19664881e-01 7.34165014e-02-5.60299551e-05    3
 2.31373796e-08-3.99759595e-12-1.71781508e+04 2.75475609e+01                   4
NC5-QOOH                C   5H  11O   2     G    300.00   3500.00 1300.00      1
 1.36538194e+01 3.77860020e-02-1.75151081e-05 3.90394425e-09-3.41708560e-13    2
-1.43879859e+04-3.94678820e+01-5.74283056e-01 8.15647789e-02-6.80290814e-05    3
 2.98085460e-08-5.32336273e-12-1.06886793e+04 3.29074336e+01                   4
NC5-OOQOOH              C   5H  11O   4     G    300.00   3500.00 1270.00      1
 1.54638476e+01 4.30531975e-02-2.04284728e-05 4.63174721e-09-4.10271992e-13    2
-3.17413365e+04-4.31406916e+01 1.43265567e+00 8.72459280e-02-7.26246112e-05    3
 3.20312949e-08-5.80388375e-12-2.81774138e+04 2.79053907e+01                   4
C4H6O2                  C   4H   6O   2     G    300.00   3500.00 1800.00      1
 7.01919581e+00 2.89919962e-02-1.39811163e-05 3.22750474e-09-2.90888809e-13    2
-4.36055710e+04-7.47846941e+00 9.15158242e-01 4.25565241e-02-2.52848896e-05    3
 7.41408744e-09-8.72358628e-13-4.14081175e+04 2.55578553e+01                   4
C4H8O                   C   4H   8O   1     G    300.00   3500.00 1800.00      1
 1.12815996e+01 2.48463701e-02-1.13234700e-05 2.47069946e-09-2.12413507e-13    2
-2.03756688e+04-3.84267373e+01-2.94845122e+00 5.64687053e-02-3.76754160e-05    3
 1.22306795e-08-1.56796629e-12-1.52528505e+04 3.85892666e+01                   4
C5H8O                   C   5H   8O   1     G    300.00   3500.00 1330.00      1
 6.70800689e+00 3.65243774e-02-1.77765821e-05 4.15639147e-09-3.79163308e-13    2
-5.52771783e+03-9.67918423e+00-5.12640161e+00 7.21165835e-02-5.79181679e-05    3
 2.42774871e-08-4.16132414e-12-2.37976516e+03 5.07899200e+01                   4
NC3H7OH                 C   3H   8O   1     G    300.00   3500.00 1800.00      1
 1.10496319e+01 1.81260731e-02-6.48607610e-06 1.10352513e-09-7.45033698e-14    2
-3.64580965e+04-3.27312856e+01-2.51644448e-01 4.32400205e-02-2.74143656e-05    3
 8.85474347e-09-1.15106147e-12-3.23896370e+04 2.84335795e+01                   4
CH3CHCH2OH              C   3H   7O   1     G    300.00   3500.00 1800.00      1
 7.63374756e+00 2.08880310e-02-8.76974163e-06 1.80199756e-09-1.48384024e-13    2
-1.08851839e+04-1.05293244e+01 2.18301336e+00 3.30007737e-02-1.88636939e-05    3
 5.54049839e-09-6.67620249e-13-8.92291955e+03 1.89711862e+01                   4
CH3CH2CHOH              C   3H   7O   1     G    300.00   3500.00 1800.00      1
 1.06992300e+01 1.62004106e-02-6.03307514e-06 1.08996004e-09-7.93898637e-14    2
-1.44167384e+04-2.94436050e+01 9.48802516e-01 3.78680272e-02-2.40894223e-05    3
 7.77749601e-09-1.00821430e-12-1.09065845e+04 2.33277424e+01                   4
CH2CH2CH2OH             C   3H   7O   1     G    300.00   3500.00 1800.00      1
 1.10024651e+01 1.50905454e-02-5.07771786e-06 7.82747262e-10-4.56159151e-14    2
-1.15495011e+04-2.90815232e+01 2.77594410e-01 3.89235914e-02-2.49385895e-05    3
 8.13862564e-09-1.06726569e-12-7.68854770e+03 2.89637142e+01                   4
CH3CH2CH2O              C   3H   7O   1     G    300.00   3500.00 1800.00      1
 6.66433268e+00 2.45624525e-02-1.14187516e-05 2.58003280e-09-2.29895788e-13    2
-7.91390086e+03-8.44862881e+00 1.62185706e+00 3.57679539e-02-2.07566695e-05    3
 6.03852088e-09-7.10241355e-13-6.09860964e+03 1.88423012e+01                   4
IC3H7OH                 C   3H   8O   1     G    300.00   3500.00 1490.00      1
 1.02736687e+01 1.89903342e-02-6.50928762e-06 9.85863990e-10-5.35101895e-14    2
-3.77812744e+04-2.92304676e+01-1.25951086e+00 4.99518902e-02-3.76786393e-05    3
 1.49318826e-08-2.39344620e-12-3.43443869e+04 3.10096138e+01                   4
CH2CHOHCH3              C   3H   7O   1     G    300.00   3500.00 1380.00      1
 6.32694430e+00 2.38762490e-02-1.07376178e-05 2.33737032e-09-2.01069469e-13    2
-1.14217376e+04-3.95690498e+00 6.40756936e-01 4.03579515e-02-2.86525118e-05    3
 1.09919085e-08-1.76892059e-12-9.85234986e+03 2.53070892e+01                   4
CH3COHCH3               C   3H   7O   1     G    300.00   3500.00 1270.00      1
 6.71652579e+00 2.35306498e-02-1.06144747e-05 2.31761627e-09-1.99886320e-13    2
-1.44175086e+04-7.90476331e+00 1.21649821e+00 4.08535713e-02-3.10746182e-05    3
 1.30578491e-08-2.31410538e-12-1.30205016e+04 1.99442900e+01                   4
C3H7CHO                 C   4H   8O   1     G    300.00   3500.00  700.00      1
-9.77279407e-01 5.24983746e-02-3.09762337e-05 8.32680249e-09-8.38156518e-13    2
-2.70767712e+04 3.27194911e+01 3.71554479e+00 2.56822364e-02 2.64869197e-05    3
-4.64000103e-08 1.87071338e-11-2.77337665e+04 1.17531399e+01                   4
RALD4X                  C   4H   7O   1     G    300.00   3500.00 1140.00      1
-3.84911251e+00 5.11968669e-02-2.73583537e-05 6.64027831e-09-6.13455715e-13    2
-5.69209146e+03 4.92440537e+01 6.06312506e+00 1.64170860e-02 1.84045160e-05    3
-2.01216338e-08 5.25538465e-12-7.95208163e+03 1.24454033e-01                   4
C3H5CHO                 C   4H   6O   1     G    300.00   3500.00 1610.00      1
 9.36564259e+00 1.99394689e-02-8.24714277e-06 1.63840913e-09-1.29181894e-13    2
-1.44293663e+04-2.07054000e+01 2.40474771e-01 4.26106933e-02-2.93694015e-05    3
 1.03846860e-08-1.48729943e-12-1.14910622e+04 2.76639767e+01                   4
IC3H5CHO                C   4H   6O   1     G    300.00   3500.00 1370.00      1
 8.96605760e+00 2.20962385e-02-1.00901145e-05 2.22139279e-09-1.91792264e-13    2
-1.79920102e+04-2.11939239e+01 6.92941976e-01 4.62513206e-02-3.65372847e-05    3
 1.50910620e-08-2.54027204e-12-1.57251765e+04 2.13235423e+01                   4
NC4H7OH                 C   4H   8O   1     G    300.00   3500.00 1260.00      1
 9.47752943e+00 2.59932961e-02-1.14395843e-05 2.45196196e-09-2.08596763e-13    2
-2.58308658e+04-2.26233180e+01-1.20059161e+00 5.98920930e-02-5.17952949e-05    3
 2.38041898e-08-4.44514991e-12-2.31399793e+04 3.13602824e+01                   4
IC4H7OH                 C   4H   8O   1     G    300.00   3500.00 1800.00      1
 1.15391986e+01 2.16392182e-02-8.55965721e-06 1.65851647e-09-1.29717162e-13    2
-2.50645509e+04-3.36074037e+01 1.41746535e+00 4.41319587e-02-2.73036076e-05    3
 8.60072033e-09-1.09391214e-12-2.14207270e+04 2.11735281e+01                   4
IC3H7CHO                C   4H   8O   1     G    300.00   3500.00 1800.00      1
 1.25375038e+01 2.06759832e-02-7.90606663e-06 1.44761601e-09-1.05776578e-13    2
-3.22363635e+04-4.10505202e+01-3.44732114e-01 4.93031741e-02-3.17620591e-05    3
 1.02831688e-08-1.33293668e-12-2.75987585e+04 2.86708279e+01                   4
RIBALDB                 C   4H   7O   1     G    300.00   3500.00 1090.00      1
 7.80130143e+00 2.08311674e-02-4.31906593e-06-1.13870083e-10 8.81387266e-14    2
-1.58031223e+03-1.28298252e+01-1.99174484e+00 5.67689519e-02-5.37747327e-05    3
 3.01342441e-08-6.84950215e-12 5.54571859e+02 3.52599043e+01                   4
RIBALDG                 C   4H   7O   1     G    300.00   3500.00 1050.00      1
 9.00440173e+00 1.88029635e-02-3.43463806e-06-2.58096325e-10 9.53220855e-14    2
-4.96767967e+03-1.61872934e+01-3.42297331e+00 6.61453446e-02-7.10666111e-05    3
 4.26828389e-08-1.01287101e-11-2.35793091e+03 4.43739411e+01                   4
N1C4H9OH                C   4H  10O   1     G    300.00   3500.00 1800.00      1
 1.48230798e+01 2.16832754e-02-7.46704085e-06 1.19388940e-09-7.36745676e-14    2
-4.08306213e+04-5.15940698e+01-4.78997489e-01 5.56878916e-02-3.58042210e-05    3
 1.16891413e-08-1.53134844e-12-3.53218735e+04 3.12239645e+01                   4
CH3CH2CHCH2OH           C   4H   9O   1     G    300.00   3500.00 1800.00      1
 1.13530982e+01 2.45578872e-02-9.82948618e-06 1.91527532e-09-1.49940483e-13    2
-1.52382167e+04-2.90980437e+01 1.95582522e+00 4.54407161e-02-2.72318436e-05    3
 8.36059288e-09-1.04512348e-12-1.18551985e+04 2.17619582e+01                   4
CH2CH2CH2CH2OH          C   4H   9O   1     G    300.00   3500.00 1790.00      1
 1.44669850e+01 1.91857603e-02-6.39892959e-06 9.65852776e-10-5.40086293e-14    2
-1.57844512e+04-4.62017057e+01 4.01250150e-02 5.14245536e-02-3.34146782e-05    3
 1.10275841e-08-1.45927837e-12-1.06196353e+04 3.17990977e+01                   4
CH3CH2CH2CH2O           C   4H   9O   1     G    300.00   3500.00 1800.00      1
 9.76394270e+00 2.97115921e-02-1.36105451e-05 3.01462692e-09-2.63554924e-13    2
-1.20864790e+04-2.37714276e+01 1.13482603e+00 4.88874069e-02-2.95903908e-05    3
 8.93308828e-09-1.08556345e-12-8.97999699e+03 2.29311520e+01                   4
CH3CH2CH2CHOH           C   4H   9O   1     G    300.00   3500.00 1800.00      1
 1.45806677e+01 1.95400847e-02-6.85981976e-06 1.13500508e-09-7.38190524e-14    2
-1.88304378e+04-4.88995705e+01 7.07705507e-01 5.03688897e-02-3.25504906e-05    3
 1.06500683e-08-1.39535562e-12-1.38361714e+04 2.61837951e+01                   4
CH3CHCH2CH2OH           C   4H   9O   1     G    300.00   3500.00 1800.00      1
 1.10474004e+01 2.49495870e-02-1.02454957e-05 2.07975625e-09-1.70767943e-13    2
-1.60937900e+04-2.75546799e+01-8.85955889e-02 4.96962447e-02-3.08677104e-05    3
 9.71761356e-09-1.23158146e-12-1.20848314e+04 3.27156533e+01                   4
N2C4H9OH                C   4H  10O   1     G    300.00   3500.00 1800.00      1
 1.39850075e+01 2.35768220e-02-8.73106105e-06 1.51546162e-09-1.02847459e-13    2
-4.24053999e+04-4.83702850e+01 1.11912947e-01 5.44059211e-02-3.44219770e-05    3
 1.10306157e-08-1.42439663e-12-3.74110858e+04 2.67137971e+01                   4
CH2CH2CHOHCH3           C   4H   9O   1     G    300.00   3500.00 1800.00      1
 1.39333095e+01 2.07599768e-02-7.56097164e-06 1.27900113e-09-8.37238499e-14    2
-1.74897435e+04-4.46134901e+01 9.11733055e-01 4.96968134e-02-3.16750021e-05    3
 1.02101235e-08-1.32415752e-12-1.28019760e+04 2.58619981e+01                   4
CH3CH2CHOHCH2           C   4H   9O   1     G    300.00   3500.00 1800.00      1
 1.39333095e+01 2.07599768e-02-7.56097164e-06 1.27900113e-09-8.37238499e-14    2
-1.74897435e+04-4.46134901e+01 9.11733055e-01 4.96968134e-02-3.16750021e-05    3
 1.02101235e-08-1.32415752e-12-1.28019760e+04 2.58619981e+01                   4
CH3CHCHOHCH3            C   4H   9O   1     G    300.00   3500.00 1800.00      1
 1.11524016e+01 2.52912378e-02-1.05179486e-05 2.12392651e-09-1.71553011e-13    2
-1.78095410e+04-2.94209720e+01 6.76902372e-01 4.85701251e-02-2.99170213e-05    3
 9.30876824e-09-1.16944770e-12-1.40383613e+04 2.72746153e+01                   4
CH3CH2COHCH3            C   4H   9O   1     G    300.00   3500.00 1430.00      1
 8.72382272e+00 3.04342830e-02-1.39185549e-05 3.06043861e-09-2.64689230e-13    2
-1.80661273e+04-1.71435098e+01 1.27395834e+00 5.12730645e-02-3.57774166e-05    3
 1.32510501e-08-2.04626467e-12-1.59354661e+04 2.14624055e+01                   4
TC4H9OH                 C   4H  10O   1     G    300.00   3500.00 1440.00      1
 9.08150387e+00 3.22201837e-02-1.41979352e-05 3.03249263e-09-2.56658356e-13    2
-4.23917231e+04-2.36263218e+01-6.99999563e-01 5.93910266e-02-4.25008966e-05    3
 1.61357155e-08-2.53152343e-12-3.95746501e+04 2.71305359e+01                   4
RTC4H8OH                C   4H   9O   1     G    300.00   3500.00 1380.00      1
 8.66823484e+00 3.01271731e-02-1.35256253e-05 2.94117291e-09-2.52822189e-13    2
-1.73478965e+04-1.68023720e+01 1.39901310e-03 5.52484364e-02-4.08313463e-05    3
 1.61323424e-08-2.64252681e-12-1.49558499e+04 2.78015457e+01                   4
IC4H9OH                 C   4H  10O   1     G    300.00   3500.00 1800.00      1
 1.44537517e+01 2.20810695e-02-7.57959310e-06 1.19533670e-09-7.16167606e-14    2
-4.15822810e+04-5.13315495e+01-5.45479447e-01 5.54126942e-02-3.53559470e-05    3
 1.14828752e-08-1.50044155e-12-3.61825578e+04 2.98474183e+01                   4
CH3CHCH3CHOH            C   4H   9O   1     G    300.00   3500.00 1450.00      1
 8.91411879e+00 2.94184843e-02-1.30488503e-05 2.81020956e-09-2.39749810e-13    2
-1.71145335e+04-1.85255698e+01 6.16106328e-01 5.23095531e-02-3.67292664e-05    3
 1.36977572e-08-2.11691319e-12-1.47081099e+04 2.45907827e+01                   4
CH3CCH2OHCH3            C   4H   9O   1     G    300.00   3500.00  700.00      1
 2.02076660e+00 4.09903684e-02-2.06486867e-05 5.00507650e-09-4.71523454e-13    2
-1.40718373e+04 2.15880988e+01 3.53447956e+00 3.23405800e-02-2.11342588e-06    3
-1.26475529e-08 5.83298703e-12-1.42837571e+04 1.48252122e+01                   4
CH2CHCH2OHCH3           C   4H   9O   1     G    300.00   3500.00 1780.00      1
 1.38129919e+01 2.02819032e-02-7.03372780e-06 1.12439860e-09-6.86002895e-14    2
-1.64045579e+04-4.42517079e+01 2.32452600e-01 5.07999690e-02-3.27511989e-05    3
 1.07564103e-08-1.42141092e-12-1.15698860e+04 2.90972641e+01                   4
MEK                     C   4H   8O   1     G    300.00   3500.00 1800.00      1
 1.00996674e+01 2.22850926e-02-8.24112797e-06 1.42760366e-09-9.77654879e-14    2
-3.40270944e+04-2.55002808e+01 1.67138626e+00 4.10146063e-02-2.38490560e-05    3
 7.20831776e-09-9.00642447e-13-3.09929132e+04 2.01153350e+01                   4
C5H9OH                  C   5H  10O   1     G    300.00   3500.00 1210.00      1
 1.31847853e+01 3.05720306e-02-1.32292735e-05 2.77400243e-09-2.30719149e-13    2
-2.99739271e+04-4.19054228e+01-3.87325759e+00 8.69622549e-02-8.31345102e-05    3
 4.12892844e-08-8.18842203e-12-2.58458807e+04 4.36413837e+01                   4
C4H9CHO                 C   5H  10O   1     G    300.00   3500.00  760.00      1
-1.78433184e+00 6.31204388e-02-3.60836199e-05 9.48321924e-09-9.39522549e-13    2
-2.97113508e+04 3.92478714e+01 5.53299033e+00 2.46082168e-02 3.99273445e-05    3
-5.71930654e-08 2.09934658e-11-3.08235838e+04 5.95416457e+00                   4
IC5H9OH                 C   5H  10O   1     G    300.00   3500.00 1340.00      1
 1.04339676e+01 3.43709884e-02-1.53823526e-05 3.33540372e-09-2.86051918e-13    2
-3.01866098e+04-2.68956309e+01-1.89607142e+00 7.11770751e-02-5.65831958e-05    3
 2.38333357e-08-4.11029295e-12-2.68821593e+04 3.61983077e+01                   4
IC4H9CHO                C   5H  10O   1     G    300.00   3500.00 1800.00      1
 1.47934378e+01 2.65660103e-02-1.04284281e-05 1.98344196e-09-1.51387846e-13    2
-3.60342983e+04-5.12505581e+01 7.73443177e-01 5.77215539e-02-3.63913811e-05    3
 1.15993505e-08-1.48693069e-12-3.09871002e+04 2.46285774e+01                   4
RALD5X                  C   5H   9O   1     G    300.00   3500.00  750.00      1
-3.04813122e-01 5.67977503e-02-3.24057644e-05 8.50471990e-09-8.41763295e-13    2
-5.21420509e+03 3.41933262e+01 6.22525357e+00 2.19707280e-02 3.72482804e-05    3
-5.34099865e-08 1.97964722e-11-6.19371509e+03 4.56811230e+00                   4
ALDC6                   C   6H  12O   1     G    300.00   3500.00 1800.00      1
 1.43376050e+01 3.78182965e-02-1.64821906e-05 3.50929997e-09-2.98005833e-13    2
-3.75955824e+04-4.53859600e+01 1.31726275e+00 6.67523904e-02-4.05939354e-05    3
 1.24395759e-08-1.53832193e-12-3.29082592e+04 2.50828483e+01                   4
RALD6X                  C   6H  11O   1     G    300.00   3500.00 1160.00      1
 5.47459470e-01 6.16901246e-02-2.98352974e-05 6.64392083e-09-5.73135815e-13    2
-1.27523068e+04 2.98980226e+01 4.05975345e+00 4.95787661e-02-1.41740579e-05    3
-2.35679152e-09 1.36667288e-12-1.35671590e+04 1.24319397e+01                   4
C5H11OH                 C   5H  12O   1     G    300.00   3500.00 1800.00      1
 1.84921366e+01 2.54355952e-02-8.57802272e-06 1.32118635e-09-7.66433346e-14    2
-4.51605186e+04-6.98750288e+01-6.77485013e-01 6.80347542e-02-4.40773219e-05    3
 1.44690750e-08-1.90273897e-12-3.82594548e+04 3.38749622e+01                   4
RPENT1OHA               C   5H  11O   1     G    300.00   3500.00 1800.00      1
 1.84065773e+01 2.29900185e-02-7.76357329e-06 1.20244128e-09-7.05741185e-14    2
-2.32226149e+04-6.80495353e+01 4.75636951e-01 6.28365526e-02-4.09690184e-05    3
 1.35007543e-08-1.77867315e-12-1.67674764e+04 2.89964546e+01                   4
RPENT1OHB               C   5H  11O   1     G    300.00   3500.00 1800.00      1
 1.50707231e+01 2.82315427e-02-1.08918053e-05 2.02927093e-09-1.51568857e-13    2
-1.95906718e+04-4.76575366e+01 1.72826109e+00 5.78814583e-02-3.56000684e-05    3
 1.11804795e-08-1.42257004e-12-1.47873854e+04 2.45546514e+01                   4
IC5H11OH                C   5H  12O   1     G    300.00   3500.00 1800.00      1
 1.75261800e+01 2.67328515e-02-9.21962742e-06 1.46158882e-09-8.81568439e-14    2
-4.58408793e+04-6.62686894e+01-6.91392019e-01 6.72163448e-02-4.29558718e-05    3
 1.39564942e-08-1.82356036e-12-3.92825534e+04 3.23286106e+01                   4
RIPENTOHA               C   5H  11O   1     G    300.00   3500.00 1620.00      1
 1.36179105e+01 3.09491059e-02-1.25439310e-05 2.45214936e-09-1.90908871e-13    2
-2.20274849e+04-4.25086987e+01 6.58084780e-01 6.29486755e-02-4.21731621e-05    3
 1.46452486e-08-2.07255998e-12-1.78285014e+04 2.62671274e+01                   4
RIPENTOHB               C   5H  11O   1     G    300.00   3500.00 1800.00      1
 1.43827445e+01 2.99341363e-02-1.24371812e-05 2.55513031e-09-2.11814101e-13    2
-2.12442482e+04-4.60019499e+01-6.44588846e-01 6.33282104e-02-4.02655763e-05    3
 1.28619433e-08-1.64331591e-12-1.58344082e+04 3.53291130e+01                   4
ESAN1OH                 C   6H  14O   1     G    300.00   3500.00 1800.00      1
 2.78613474e+01 1.77437818e-02-2.99502852e-06 1.18974668e-11 2.84572872e-14    2
-5.19282550e+04-1.19896980e+02-1.83303781e+00 8.37313045e-02-5.79846308e-05    3
 2.03784168e-08-2.80022596e-12-4.12382763e+04 4.08152273e+01                   4
RESAN1OHA               C   6H  13O   1     G    300.00   3500.00 1800.00      1
 2.84298178e+01 1.33218304e-02-9.68178066e-07-3.32583082e-10 4.90833295e-14    2
-3.02913834e+04-1.20327849e+02-1.87679570e-01 7.69162690e-02-5.39635435e-05    3
 1.92953301e-08-2.67701572e-12-1.99890844e+04 3.45560167e+01                   4
RESAN1OHB               C   6H  13O   1     G    300.00   3500.00 1800.00      1
 2.97416428e+01 1.08284395e-02 6.26458140e-07-7.76125692e-10 9.43842404e-14    2
-2.87904782e+04-1.27477419e+02-8.09485399e-02 7.71008646e-02-5.46005628e-05    3
 1.96783265e-08-2.74651190e-12-1.80543453e+04 3.39286664e+01                   4
NC5H12                  C   5H  12          G    300.00   3500.00 1800.00      1
 2.12559082e+01 1.49866375e-02-1.56738310e-06-4.84518439e-10 9.00436513e-14    2
-2.80668702e+04-9.05497671e+01-1.97000865e+00 6.65997861e-02-4.45783403e-05    3
 1.54454657e-08-2.12245414e-12-1.97055401e+04 3.51537401e+01                   4
NC5H11                  C   5H  11          G    300.00   3500.00 1800.00      1
 6.93193785e+00 3.75440987e-02-1.65478566e-05 3.53633643e-09-2.99976701e-13    2
-1.73087074e+03-8.88710671e+00-3.57520449e+00 6.08933039e-02-3.60055276e-05    3
 1.07428812e-08-1.30088570e-12 2.05170050e+03 4.79797395e+01                   4
NEOC5H12                C   5H  12          G    300.00   3500.00 1700.00      1
 1.58220811e+01 2.73824077e-02-1.01392581e-05 1.77707009e-09-1.22756971e-13    2
-2.85197010e+04-6.62488521e+01-2.62463459e+00 7.07864445e-02-4.84369376e-05    3
 1.67957680e-08-2.33138901e-12-2.22478177e+04 3.25342362e+01                   4
NEOC5H11                C   5H  11          G    300.00   3500.00 1670.00      1
 1.43276289e+01 2.66845577e-02-1.02158264e-05 1.86929104e-09-1.35803312e-13    2
-2.94216421e+03-5.15145769e+01-1.29689709e+00 6.41085720e-02-4.38302105e-05    3
 1.52882069e-08-2.14462305e-12 2.27642747e+03 3.18773552e+01                   4
NC5H10                  C   5H  10          G    300.00   3500.00 1800.00      1
 1.11929736e+01 2.82582223e-02-1.13863841e-05 2.22526491e-09-1.74280993e-13    2
-1.02483443e+04-3.39253533e+01-6.89551965e-01 5.46638348e-02-3.33910611e-05    3
 1.03751453e-08-1.30620882e-12-5.97063504e+03 3.03853541e+01                   4
NC5H9-3                 C   5H   9          G    300.00   3500.00 1800.00      1
 9.88287390e+00 2.86275350e-02-1.23662428e-05 2.58308509e-09-2.14520963e-13    2
 7.14211639e+03-2.81379758e+01-9.61360662e-01 5.27258341e-02-3.24481586e-05    3
 1.00208317e-08-1.24754133e-12 1.10460408e+04 3.05532839e+01                   4
B1M2                    C   5H  10          G    300.00   3500.00 1800.00      1
 1.21299340e+01 2.65376145e-02-1.02995525e-05 1.93064538e-09-1.45051208e-13    2
-1.11266091e+04-3.96207198e+01-6.39002025e-01 5.49130280e-02-3.39457304e-05    3
 1.06884890e-08-1.36141838e-12-6.52979211e+03 2.94874259e+01                   4
B1M3                    C   5H  10          G    300.00   3500.00 1800.00      1
 1.31681365e+01 2.49963287e-02-9.30063098e-06 1.64277853e-09-1.14892348e-13    2
-1.09953810e+04-4.60629131e+01-8.44094903e-01 5.61346208e-02-3.52492077e-05    3
 1.12533625e-08-1.44969568e-12-5.95097767e+03 2.97742066e+01                   4
B2M2                    C   5H  10          G    300.00   3500.00 1800.00      1
 9.73411699e+00 3.08235227e-02-1.30972997e-05 2.71635425e-09-2.25270435e-13    2
-1.14704814e+04-2.74877025e+01 1.14407401e-01 5.22006552e-02-3.09115767e-05    3
 9.31423462e-09-1.14164271e-12-8.00738598e+03 2.45761726e+01                   4
CYC5H8                  C   5H   8          G    300.00   3500.00 1460.00      1
 8.43099916e+00 2.71082714e-02-1.07932861e-05 1.95387665e-09-1.31111174e-13    2
-1.09862538e+03-2.37608448e+01-6.56863981e+00 6.82031726e-02-5.30140751e-05    3
 2.12327757e-08-3.43229252e-12 3.28126920e+03 5.42801525e+01                   4
C5H7                    C   5H   7          G    300.00   3500.00 1430.00      1
 7.72404526e+00 2.56072196e-02-8.76350315e-06 8.66193956e-10 3.30416653e-14    2
 2.30808142e+04-1.69352935e+01 2.31765046e-01 4.65646468e-02-3.07468184e-05    3
 1.11148258e-08-1.75867718e-12 2.52236063e+04 2.18904247e+01                   4
LC5H8                   C   5H   8          G    300.00   3500.00 1430.00      1
 8.95829160e+00 2.51033002e-02-8.43679233e-06 8.19905618e-10 3.11426514e-14    2
 4.67953300e+03-2.40439629e+01 1.19183501e+00 4.68276543e-02-3.12245763e-05    3
 1.14435811e-08-1.82614328e-12 6.90073958e+03 1.62025638e+01                   4
DIALLYL                 C   6H  10          G    300.00   3500.00 1670.00      1
 1.46885479e+01 2.58341295e-02-9.34005191e-06 1.60362032e-09-1.08722036e-13    2
 2.72208305e+03-5.11904321e+01-8.93391062e-01 6.31561390e-02-4.28628150e-05    3
 1.49859609e-08-2.11206643e-12 7.92645066e+03 3.19742028e+01                   4
RC6H9A                  C   6H   9          G    300.00   3500.00 1310.00      1
 1.02179198e+01 3.31131696e-02-1.50182300e-05 3.28859653e-09-2.83959224e-13    2
 2.30740211e+04-2.53806643e+01-2.61882183e+00 7.23093274e-02-5.98993266e-05    3
 2.61288493e-08-4.64278609e-12 2.64372474e+04 4.00154625e+01                   4
CYC6H8                  C   6H   8          G    300.00   3500.00 1490.00      1
 8.66772261e+00 3.45074855e-02-1.63846780e-05 3.69260974e-09-3.24421025e-13    2
 5.74022138e+03-2.73566208e+01-6.91358136e+00 7.63364895e-02-5.84944135e-05    3
 2.25336547e-08-3.48567018e-12 1.03834500e+04 5.40276160e+01                   4
CYC6H10                 C   6H  10          G    300.00   3500.00 1800.00      1
 1.51624858e+01 2.76360017e-02-1.05259858e-05 1.89586361e-09-1.35054774e-13    2
-9.29985244e+03-6.25064559e+01-6.01517655e+00 7.46974737e-02-4.97438791e-05    3
 1.64210093e-08-2.15243611e-12-1.67589399e+03 5.21114707e+01                   4
RCYC6H9                 C   6H   9          G    300.00   3500.00 1800.00      1
 1.41670463e+01 2.75651338e-02-1.13337615e-05 2.23021652e-09-1.74683445e-13    2
 7.93866332e+03-5.85441979e+01-6.48639356e+00 7.34616669e-02-4.95808724e-05    3
 1.63958131e-08-2.14212742e-12 1.53739017e+04 5.32365273e+01                   4
CYC6H12                 C   6H  12          G    300.00   3500.00 1800.00      1
 1.12578097e+01 4.34354098e-02-2.02455774e-05 4.54245292e-09-4.01195170e-13    2
-2.30439963e+04-4.47863376e+01-9.43363126e+00 8.94163897e-02-5.85630607e-05    3
 1.87341134e-08-2.37225913e-12-1.55950776e+04 6.72000574e+01                   4
CYC6H11                 C   6H  11          G    300.00   3500.00 1800.00      1
 1.12879191e+01 3.94798364e-02-1.80474738e-05 3.97976998e-09-3.47933572e-13    2
 4.69934404e+02-4.15743644e+01-9.20200373e+00 8.50129981e-02-5.59917752e-05    3
 1.80332150e-08-2.29980093e-12 7.84630661e+03 6.93213721e+01                   4
NC6H12                  C   6H  12          G    300.00   3500.00 1780.00      1
 2.80951655e+01 5.24635940e-03 6.43208140e-06-3.19131390e-09 4.01093698e-13    2
-1.79767847e+04-1.24497292e+02-1.85358315e+00 7.25469181e-02-5.02818725e-05    3
 1.80498674e-08-2.58221828e-12-7.31503024e+03 3.72569567e+01                   4
NC7H16                  C   7H  16          G    300.00   3500.00 1800.00      1
 3.10696120e+01 1.73458864e-02-4.57663866e-07-1.06280964e-09 1.59098857e-13    2
-3.76541592e+04-1.40920498e+02-2.76912812e+00 9.25430866e-02-6.31219974e-05    3
 2.21462028e-08-3.06437509e-12-2.54722127e+04 4.22218230e+01                   4
NC7H15                  C   7H  15          G    300.00   3500.00 1800.00      1
 1.58938298e+01 4.32851195e-02-1.83429598e-05 3.81524631e-09-3.18291961e-13    2
-8.33589206e+03-5.34387877e+01-1.03213606e+00 8.08983770e-02-4.96873411e-05    3
 1.54242764e-08-1.93065725e-12-2.24254435e+03 3.81680706e+01                   4
NC7H14                  C   7H  14          G    300.00   3500.00 1800.00      1
 1.82668105e+01 3.59607889e-02-1.37346402e-05 2.52229049e-09-1.85248240e-13    2
-1.87497345e+04-6.92309266e+01-1.22797310e+00 7.92825302e-02-4.98360912e-05    3
 1.58931983e-08-2.04231877e-12-1.17316124e+04 3.62789089e+01                   4
NC7H13                  C   7H  13          G    300.00   3500.00 1800.00      1
 9.88287390e+00 2.86275350e-02-1.23662428e-05 2.58308509e-09-2.14520963e-13    2
 7.14211639e+03-2.81379758e+01-9.61360662e-01 5.27258341e-02-3.24481586e-05    3
 1.00208317e-08-1.24754133e-12 1.10460408e+04 3.05532839e+01                   4
IC8H18                  C   8H  18          G    300.00   3500.00 1390.00      1
 2.06155885e+01 4.43694094e-02-1.35968858e-05 1.75327621e-09-6.83090867e-14    2
-3.76580614e+04-8.42148794e+01-5.96912082e+00 1.20872170e-01-9.61538218e-05    3
 4.13489290e-08-7.18982937e-12-3.02675122e+04 5.27954202e+01                   4
IC8H17                  C   8H  17          G    300.00   3500.00 1530.00      1
 2.65104230e+01 3.01796816e-02-5.82184988e-06 1.42085775e-11 7.60110768e-14    2
-1.80373025e+04-1.14981197e+02-3.32961207e+00 1.08192845e-01-8.23053436e-05    3
 3.33403496e-08-5.36943681e-12-8.90625182e+03 4.16697270e+01                   4
IC8H16                  C   8H  16          G    300.00   3500.00 1400.00      1
 1.88616063e+01 4.14292819e-02-1.28170543e-05 1.66806735e-09-6.58961701e-14    2
-2.24684067e+04-7.38514297e+01-5.35586582e+00 1.10622059e-01-8.69521730e-05    3
 3.69705048e-08-6.36990286e-12-1.56875145e+04 5.11323812e+01                   4
DIMEPTD                 C   7H  12          G    300.00   3500.00 1310.00      1
 1.53755546e+01 3.27318282e-02-1.05955708e-05 1.52102629e-09-7.69415904e-14    2
-6.19682930e+03-5.37226047e+01-1.29247814e+00 8.36265847e-02-6.88720095e-05    3
 3.11782470e-08-5.73671653e-12-1.82980473e+03 3.11918394e+01                   4
C7H8                    C   7H   8          G    200.00   3500.00 1740.00      1
 1.92535108e+01 1.64137602e-02-3.61135948e-06 2.27424890e-11 5.04456794e-14    2
-3.67626229e+03-8.27561068e+01-4.42382865e+00 7.08444256e-02-5.05343469e-05    3
 1.80008986e-08-2.53262272e-12 4.56345183e+03 4.45878951e+01                   4
C6H5OH                  C   6H   6O   1     G    300.00   3500.00 1330.00      1
 1.39867713e+01 2.02277643e-02-7.36599497e-06 1.21196287e-09-7.46105009e-14    2
-1.80542263e+04-5.08485812e+01-5.47325436e+00 7.87541571e-02-7.33732049e-05    3
 3.42982837e-08-6.29384373e-12-1.28778595e+04 4.85843830e+01                   4
C6H5CHO                 C   7H   6O   1     G    200.00   3500.00 1630.00      1
 2.06104936e+01 1.34209230e-02-2.83635978e-06-5.48103780e-11 5.23167108e-14    2
-1.43315560e+04-8.70895599e+01-3.50845143e+00 7.26085180e-02-5.73034718e-05    3
 2.22221271e-08-3.36439149e-12-6.46877992e+03 4.10544422e+01                   4
C6H5CO                  C   7H   5O   1     G    300.00   3500.00 1470.00      1
 1.31799087e+01 2.42895707e-02-1.09067387e-05 2.35371847e-09-2.00195165e-13    2
 5.86598787e+03-4.37756649e+01-1.56203256e+00 6.44036967e-02-5.18395203e-05    3
 2.09173383e-08-3.35727336e-12 1.02001186e+04 3.30251959e+01                   4
C7H7                    C   7H   7          G    200.00   3500.00 1600.00      1
 1.77148781e+01 1.72901839e-02-4.74309316e-06 3.88421745e-10 1.27959347e-14    2
 1.68881058e+04-7.24712964e+01-3.23806381e+00 6.96725387e-02-5.38515508e-05    3
 2.08502791e-08-3.18436927e-12 2.35930472e+04 3.84624951e+01                   4
CH3C6H4                 C   7H   7          G    200.00   3500.00 1730.00      1
 1.83842182e+01 1.52647348e-02-3.43004339e-06 5.73661650e-11 4.21798063e-14    2
 2.84624024e+04-7.44700925e+01-2.82564598e+00 6.43048832e-02-4.59504033e-05    3
 1.64428613e-08-2.32566631e-12 3.58010154e+04 3.94808224e+01                   4
C6H5O                   H   5C   6O   1     G    100.00   3500.00 1800.00      1
 1.20320192e+01 2.29423311e-02-1.10171059e-05 2.53057377e-09-2.25735901e-13    2
 2.17286268e+02-4.10084349e+01 4.06305309e-01 4.87772509e-02-3.25462057e-05    3
 1.05043144e-08-1.33319988e-12 4.40254327e+03 2.19123540e+01                   4
BENZYNE                 C   6H   4          G    300.00   3500.00 1400.00      1
 1.09465819e+01 1.50373245e-02-5.27844957e-06 8.14607575e-10-4.49073360e-14    2
 5.03301418e+04-3.53782935e+01-3.73796174e+00 5.69931634e-02-5.02311341e-05    3
 2.22206478e-08-3.86741452e-12 5.44418140e+04 4.04070822e+01                   4
RCATEC                  C   6H   5O   2     G    300.00   3500.00 1140.00      1
 1.40810369e+01 2.16036557e-02-9.34848721e-06 1.81734387e-09-1.31737733e-13    2
-2.57458618e+04-4.55416676e+01-4.82568618e+00 8.79430349e-02-9.66371440e-05    3
 5.28633420e-08-1.13260356e-11-2.14351289e+04 4.81496572e+01                   4
C6H4O2                  C   6H   4O   2     G    300.00   3500.00 1410.00      1
 1.74929578e+01 1.29021286e-02-2.02976640e-06-3.72417853e-10 8.59745736e-14    2
-2.22100459e+04-6.49015838e+01-5.23446579e+00 7.73770890e-02-7.06201498e-05    3
 3.20580235e-08-5.66410368e-12-1.58009124e+04 5.25540058e+01                   4
CYC5H4O                 C   5H   4O   1     G    300.00   3500.00 1260.00      1
 6.34459580e+00 2.39841575e-02-8.32755386e-06 8.47127646e-10 2.86249491e-14    2
 3.08659308e+03-9.73181560e+00-5.14379340e+00 6.04552343e-02-5.17455025e-05    3
 2.38195872e-08-4.52940274e-12 5.98166715e+03 4.83481228e+01                   4
C7H7O2                  C   7H   7O   2     G    300.00   3500.00 1420.00      1
 1.76964624e+01 2.58808958e-02-1.00755993e-05 1.78285132e-09-1.17592477e-13    2
 6.43630911e+03-6.45881471e+01-4.45172572e+00 8.82701582e-02-7.59797497e-05    3
 3.27237670e-08-5.56493679e-12 1.27263945e+04 5.00304723e+01                   4
O2C6H4CH3               C   7H   7O   2     G    300.00   3500.00 1300.00      1
 1.57011694e+01 2.91723896e-02-1.27991927e-05 2.73382155e-09-2.31734775e-13    2
 5.63564260e+03-5.46747931e+01-5.21645096e+00 9.35342985e-02-8.70629336e-05    3
 4.08177913e-08-7.55557510e-12 1.10742239e+04 5.17286697e+01                   4
OC6H4CH2                C   7H   6O   1     G    300.00   3500.00 1390.00      1
 1.45795344e+01 2.32519437e-02-8.58329372e-06 1.38947459e-09-7.81466970e-14    2
-5.01093188e+02-5.31869652e+01-4.82277790e+00 7.90859360e-02-6.88358034e-05    3
 3.02875608e-08-5.27564421e-12 4.89274964e+03 4.68072303e+01                   4
C6H5CH2O                C   7H   7O   1     G    300.00   3500.00 1650.00      1
 1.54569227e+01 2.51288522e-02-9.88344275e-06 1.85206220e-09-1.37473827e-13    2
 6.00712849e+03-5.64457004e+01-4.49397764e+00 7.34946712e-02-5.38523691e-05    3
 1.96172850e-08-2.82917425e-12 1.25909256e+04 4.97967788e+01                   4
BZCOOH                  C   7H   8O   2     G    300.00   3500.00 1550.00      1
 1.78036107e+01 3.06807111e-02-1.34555335e-05 2.81495360e-09-2.31878498e-13    2
-1.15055065e+04-6.47324084e+01-3.42659307e+00 8.54683337e-02-6.64758135e-05    3
 2.56193751e-08-3.91001099e-12-4.92414334e+03 4.69952939e+01                   4
C6H5O2                  C   6H   5O   2     G    300.00   3500.00 1300.00      1
 1.17436568e+01 2.50264983e-02-1.11158434e-05 2.39771212e-09-2.04780348e-13    2
 1.03023085e+04-3.29345582e+01-2.98072562e+00 7.03322902e-02-6.33917571e-05    3
 2.92058730e-08-5.36019590e-12 1.41306479e+04 4.19652270e+01                   4
RBBENZ                  C  14H  13          G    300.00   3500.00 1750.00      1
 5.34298872e+01-2.73976091e-03 1.40930518e-05-5.29858386e-09 5.98002536e-13    2
 9.33192271e+03-2.64139662e+02-8.67312060e+00 1.39209971e-01-1.07578147e-04    3
 4.10523491e-08-6.02355932e-12 3.10679755e+04 7.02252758e+01                   4
STILB                   C  14H  12          G    300.00   3500.00 1470.00      1
 3.31295359e+01 3.16424147e-02-7.88066870e-06 4.81370280e-10 4.43949941e-14    2
 1.37146851e+04-1.52659599e+02-1.11031623e+01 1.52003498e-01-1.30698101e-04    3
 5.61808860e-08-9.42831176e-12 2.67190984e+04 7.77787968e+01                   4
OOC6H4OH                H   5C   6O   3     G    100.00   3500.00 1570.00      1
 2.76569225e+01 2.91346366e-04 5.46428411e-06-2.09157763e-09 2.40972768e-13    2
-1.39658758e+04-1.18517523e+02-4.81896279e-01 7.19826044e-02-6.30305484e-05    3
 2.69932769e-08-4.39037350e-12-5.13028675e+03 2.99287472e+01                   4
C6H4OH                  C   6H   5O   1     G    300.00   3500.00 1170.00      1
 1.35501563e+01 1.98692226e-02-8.43356667e-06 1.70584597e-09-1.35582641e-13    2
 1.32571078e+04-4.75538960e+01-6.19433347e+00 8.73717517e-02-9.49752706e-05    3
 5.10173582e-08-1.06722306e-11 1.78773184e+04 5.08018126e+01                   4
C7H6                    C   7H   6          G    300.00   3500.00 1290.00      1
 1.11282362e+01 2.73165807e-02-1.25329645e-05 2.76951413e-09-2.40721375e-13    2
 3.69620905e+04-3.50553513e+01-3.97785296e+00 7.41571673e-02-6.69987629e-05    3
 3.09172135e-08-5.69570188e-12 4.08594615e+04 4.16694449e+01                   4
C7H5                    C   7H   5          G    300.00   3500.00 1250.00      1
 1.21079560e+01 2.22665290e-02-9.87308079e-06 2.11666746e-09-1.79360812e-13    2
 5.15977924e+04-3.78517160e+01-2.81419579e+00 7.00174146e-02-6.71741435e-05    3
 3.26772342e-08-6.29147417e-12 5.53283304e+04 3.74688223e+01                   4
CYC5H4                  C   5H   4          G    200.00   3500.00 1310.00      1
 6.52292971e+00 1.75112092e-02-7.24525150e-06 1.36813992e-09-9.77801509e-14    2
 6.01459585e+04-1.09295493e+01-1.67820643e+00 4.25528463e-02-3.59188817e-05    3
 1.59603181e-08-2.88254699e-12 6.22946562e+04 3.08507212e+01                   4
C5H3                    C   5H   3          G    300.00   3500.00 1370.00      1
 1.06729929e+01 9.74586302e-03-3.33881730e-06 5.09387247e-10-2.86889361e-14    2
 6.39774214e+04-2.94129104e+01 3.35962353e+00 3.10987662e-02-2.67179083e-05    3
 1.18860739e-08-2.10472664e-12 6.59812846e+04 8.17219633e+00                   4
C5H2                    C   5H   2          G    300.00   3500.00 1260.00      1
 1.08586495e+01 8.25356562e-03-3.15379453e-06 5.51063161e-10-3.71272440e-14    2
 7.89908994e+04-3.35264726e+01 1.78531794e+00 3.70577929e-02-3.74445412e-05    3
 1.86943154e-08-3.63697888e-12 8.12773789e+04 1.23440607e+01                   4
C5H5O                   C   5H   5O   1     G    300.00   3500.00 1450.00      1
 1.05801390e+01 2.13128784e-02-9.63052935e-06 2.09384798e-09-1.79321203e-13    2
 1.62543411e+04-3.26154734e+01-4.01979397e+00 6.15885556e-02-5.12950230e-05    3
 2.12499370e-08-3.48209517e-12 2.04883217e+04 4.32455666e+01                   4
LC6H6                   C   6H   6          G    300.00   3500.00 1250.00      1
 1.28863876e+01 1.90072460e-02-7.30992555e-06 1.31482494e-09-9.21385778e-14    2
 3.55364843e+04-4.09021933e+01-1.05889384e+00 6.36321466e-02-6.08598063e-05    3
 2.98747613e-08-5.80412586e-12 3.90228046e+04 2.94875281e+01                   4
C6H4C2H3                C   8H   7          G    200.00   3500.00 1580.00      1
 1.99256075e+01 1.67315530e-02-4.18312961e-06 2.15370099e-10 3.07179808e-14    2
 3.89930312e+04-8.19571079e+01-3.96125911e+00 7.72046330e-02-6.15942816e-05    3
 2.44394849e-08-3.80221157e-12 4.65412811e+04 4.42096620e+01                   4
CRESOL                  C   7H   8O   1     G    300.00   3500.00 1310.00      1
 1.22673687e+01 3.34155282e-02-1.38949870e-05 2.56768165e-09-1.71519558e-13    2
-2.17187243e+04-3.95715125e+01-4.41843936e+00 8.43645604e-02-7.22335735e-05    3
 3.22565297e-08-5.83733026e-12-1.73470426e+04 4.54334870e+01                   4
RCRESOLC                C   7H   7O   1     G    300.00   3500.00 1150.00      1
 1.31541709e+01 2.50657189e-02-5.32353909e-06-2.12687604e-10 1.25840461e-13    2
-3.38086419e+03-4.22339553e+01-6.42956807e+00 9.31830718e-02-9.41722602e-05    3
 5.12938174e-08-1.10712258e-11 1.12339577e+03 5.49833260e+01                   4
RCRESOLO                C   7H   7O   1     G    300.00   3500.00 1150.00      1
 1.27824814e+01 2.40796407e-02-4.51347940e-06-4.25076353e-10 1.44988491e-13    2
-3.97704754e+03-4.00543784e+01-6.60757191e+00 9.15233043e-02-9.24834754e-05    3
 5.05720228e-08-1.09413374e-11 4.82664712e+02 5.62014117e+01                   4
C6H5CH2OH               C   7H   8O   1     G    300.00   3500.00 1450.00      1
 1.25818443e+01 2.64134519e-02-7.93799877e-06 4.38368234e-10 8.64078966e-14    2
-1.87828963e+04-3.81332334e+01-6.02884975e+00 7.77532977e-02-6.10481841e-05    3
 2.48568442e-08-4.12367417e-12-1.33857950e+04 5.85676633e+01                   4
C6H5C2H                 C   8H   6          G    200.00   3500.00 1280.00      1
 1.52608076e+01 2.33328927e-02-9.12947230e-06 1.67060897e-09-1.19620450e-13    2
 3.14643486e+04-5.61979008e+01-2.98097334e+00 8.03384582e-02-7.59328693e-05    3
 3.64640449e-08-6.91521341e-12 3.61342445e+04 3.63113150e+01                   4
C6H4C2H                 C   8H   5          G    200.00   3500.00 1410.00      1
 1.60102852e+01 1.80276839e-02-6.10631287e-06 8.89485624e-10-4.39310921e-14    2
 6.01004863e+04-5.91795508e+01-2.59308039e+00 7.08031891e-02-6.22504674e-05    3
 2.74351852e-08-4.75061541e-12 6.53466354e+04 3.69628594e+01                   4
C6H5C2H3                C   8H   8          G    200.00   3500.00 1620.00      1
 2.08689853e+01 1.76153525e-02-4.02709967e-06 7.62333198e-11 4.96213073e-14    2
 7.92336685e+03-8.97908225e+01-4.75261288e+00 8.08785579e-02-6.26041417e-05    3
 2.41820119e-08-3.67040626e-12 1.62247647e+04 4.61791070e+01                   4
C6H5C2H5                C   8H  10          G    200.00   3500.00 1660.00      1
 2.15526224e+01 2.25377527e-02-5.71678491e-06 3.25228910e-10 3.67333515e-14    2
-7.08672427e+03-9.37205827e+01-4.75947977e+00 8.59404087e-02-6.30083415e-05    3
 2.33338862e-08-3.42842587e-12 1.64889367e+03 4.65555372e+01                   4
C6H5C2H2                C   8H   7          G    200.00   3500.00 1520.00      1
 1.92541493e+01 1.80154928e-02-5.00513523e-06 4.35360010e-10 9.55509220e-15    2
 3.83998804e+04-7.81182474e+01-4.29898225e+00 7.99974179e-02-6.61715087e-05    3
 2.72627168e-08-4.40283911e-12 4.55600324e+04 4.53739369e+01                   4
C6H5CHCH3               C   8H   9          G    200.00   3500.00 1700.00      1
 2.17404159e+01 1.87953891e-02-4.10981050e-06 2.63149780e-14 6.24669644e-14    2
 1.18126541e+04-9.21825395e+01-3.04486857e+00 7.71137055e-02-5.55671485e-05    3
 2.01793745e-08-2.90508425e-12 2.02396509e+04 4.05439030e+01                   4
XYLENE                  C   8H  10          G    200.00   3500.00 1800.00      1
 2.00142025e+01 2.37296570e-02-6.76483884e-06 7.09529215e-10-1.05911395e-14    2
-8.30085767e+03-8.55893311e+01-3.92128796e+00 7.69196357e-02-5.10898211e-05    3
 1.71261893e-08-2.29068282e-12 3.15918887e+02 4.39545364e+01                   4
RXYLENE                 C   8H   9          G    200.00   3500.00 1620.00      1
 2.04972497e+01 2.14206934e-02-5.61362086e-06 3.90126528e-10 2.53125355e-14    2
 1.19614465e+04-8.71674754e+01-3.85447699e+00 8.15484138e-02-6.12874360e-05    3
 2.33011616e-08-3.51034102e-12 1.98514059e+04 4.20634392e+01                   4
INDENE                  C   9H   8          G    200.00   3500.00 1610.00      1
 2.31048443e+01 1.91297591e-02-4.53548120e-06 1.22196710e-10 5.15078704e-14    2
 8.53092089e+03-1.04304478e+02-6.87762290e+00 9.36203608e-02-7.39366630e-05    3
 2.88597461e-08-4.41084452e-12 1.81852753e+04 5.46222708e+01                   4
INDENYL                 C   9H   7          G    200.00   3500.00 1430.00      1
 2.02650248e+01 2.20602643e-02-7.28401475e-06 9.93375839e-10-4.12199483e-14    2
 2.49669757e+04-8.59379552e+01-6.82385337e+00 9.78333502e-02-8.67662727e-05    3
 3.80480416e-08-6.51930836e-12 3.27143949e+04 5.44392228e+01                   4
C10H7                   C  10H   7          G    200.00   3500.00 1490.00      1
 2.12397127e+01 2.27484190e-02-6.96640086e-06 8.04033892e-10-1.68765826e-14    2
 3.76445830e+04-9.11799918e+01-6.45168838e+00 9.70877508e-02-8.18046543e-05    3
 3.42887110e-08-5.63511100e-12 4.58966205e+04 5.34576808e+01                   4
C10H7OH                 C  10H   8O   1     G    300.00   3500.00 1730.00      1
 2.61818224e+01 2.47079229e-02-8.75472975e-06 1.41213209e-09-8.61580367e-14    2
-1.58338687e+04-1.19314317e+02-3.09194614e+00 9.23929369e-02-6.74411581e-05    3
 2.40273261e-08-3.35424965e-12-5.70514482e+03 3.79602738e+01                   4
C10H7O                  C  10H   7O   1     G    200.00   3500.00 1520.00      1
 2.51245261e+01 2.12349446e-02-5.95579175e-06 5.14900720e-10 1.27936894e-14    2
 2.27944423e+03-1.11444345e+02-6.17635896e+00 1.03605695e-01-8.72427162e-05    3
 3.61670606e-08-5.85104839e-12 1.17949133e+04 5.26703358e+01                   4
C10H6CH3                C  11H   9          G    200.00   3500.00 1530.00      1
 2.52493034e+01 2.50352394e-02-6.91797177e-06 5.80757389e-10 1.70685086e-14    2
 3.22365770e+04-1.13732286e+02-6.94188403e+00 1.09195207e-01-8.94277435e-05    3
 3.65327276e-08-5.85743643e-12 4.20870803e+04 5.52614582e+01                   4
C10H7CH2                C  11H   9          G    200.00   3500.00 1480.00      1
 2.49658354e+01 2.73321443e-02-8.56500981e-06 1.05181516e-09-3.08784850e-14    2
 2.10853669e+04-1.11434350e+02-7.41870774e+00 1.14857936e-01-9.72735830e-05    3
 4.10106319e-08-6.78067861e-12 3.06711917e+04 5.74984546e+01                   4
C10H7CHO                C  11H   8O   1     G    200.00   3500.00 1700.00      1
 3.52801173e+01 1.31180999e-02-5.97608673e-07-9.89256296e-10 1.64132767e-13    2
-1.29136404e+04-1.70276910e+02-6.53399067e+00 1.11504236e-01-8.74089056e-05    3
 3.30543895e-08-4.84228574e-12 1.30315629e+03 5.36397371e+01                   4
C10H7CH3                C  11H  10          G    200.00   3500.00 1700.00      1
 3.19556671e+01 1.89589747e-02-2.92887930e-06-5.41537998e-10 1.30075116e-13    2
-1.51641167e+03-1.52538802e+02-7.17710534e+00 1.11036086e-01-8.41733896e-05    3
 3.13190543e-08-4.55530610e-12 1.17887310e+04 5.70191587e+01                   4
CH3C10H6OH              C  11H  10O   1     G    300.00   3500.00 1800.00      1
 2.91191869e+01 2.86451308e-02-9.80098219e-06 1.51374083e-09-8.72237945e-14    2
-2.13626711e+04-1.32660114e+02-1.76841814e+00 9.72842531e-02-6.70002508e-05    3
 2.26986551e-08-3.02957300e-12-1.02431333e+04 3.45100483e+01                   4
CH3C10H6O               C  11H   9O   1     G    300.00   3500.00 1800.00      1
 2.60936624e+01 3.24954978e-02-1.30480618e-05 2.52260906e-09-1.95492396e-13    2
-2.87396993e+03-1.14905139e+02-1.85059487e+00 9.45938472e-02-6.47966864e-05    3
 2.16887663e-08-2.85745868e-12 7.18596268e+03 3.63350107e+01                   4
C12H8                   C  12H   8          G    200.00   3500.00 1570.00      1
 2.77000801e+01 2.26169409e-02-5.57154154e-06 2.34725134e-10 5.00956725e-14    2
 1.79557632e+04-1.32407942e+02-8.95027490e+00 1.15993641e-01-9.47849497e-05    3
 3.81172764e-08-5.98215771e-12 2.94639746e+04 6.09409166e+01                   4
C12H7                   C  12H   7          G    200.00   3500.00 1550.00      1
 2.72643903e+01 2.07706175e-02-5.09002113e-06 1.94274019e-10 4.95146521e-14    2
 5.03500896e+04-1.28964295e+02-8.21375630e+00 1.12327125e-01-9.36930927e-05    3
 3.83031220e-08-6.09707373e-12 6.13483151e+04 5.77457270e+01                   4
BIPHENYL                C  12H  10          G    200.00   3500.00 1620.00      1
 3.03550325e+01 2.42378629e-02-5.78855002e-06 1.73424746e-10 6.27217930e-14    2
 7.33500914e+03-1.42781766e+02-7.48580974e+00 1.17672041e-01-9.23016780e-05    3
 3.57755350e-08-5.43143103e-12 1.95954420e+04 5.80338349e+01                   4
C12H9                   C  12H   9          G    300.00   3500.00 1430.00      1
 2.37129726e+01 3.27032394e-02-1.16108738e-05 1.80515253e-09-1.00356246e-13    2
 4.00500330e+04-1.02303886e+02-9.58279780e+00 1.25838261e-01-1.09304953e-04    3
 4.73501778e-08-8.06277324e-12 4.95726233e+04 7.02380051e+01                   4
FLUORENE                C  13H  10          G    200.00   3500.00 1580.00      1
 3.04981916e+01 2.54134515e-02-6.12250971e-06 2.13473325e-10 6.26029968e-14    2
 6.42406071e+03-1.44876912e+02-9.12299946e+00 1.25720264e-01-1.01350497e-04    3
 4.03940585e-08-6.29508454e-12 1.89443571e+04 6.43961494e+01                   4
C6H5CH2C6H5             C  13H  12          G    200.00   3500.00 1730.00      1
 3.68978946e+01 2.09448951e-02-2.15140891e-06-1.01983321e-09 1.90993351e-13    2
 1.61235408e+03-1.77722051e+02-9.21937242e+00 1.27574414e-01-9.46047492e-05    3
 3.46076582e-08-4.95748807e-12 1.75689285e+04 7.00449656e+01                   4
C14H10                  C  14H  10          G    200.00   3500.00 1550.00      1
 3.33910328e+01 2.79675689e-02-7.16206047e-06 3.83005680e-10 5.29481034e-14    2
 8.53646106e+03-1.60739744e+02-9.79770356e+00 1.39422372e-01-1.15021548e-04    3
 4.67741830e-08-7.42949985e-12 2.19249693e+04 6.65486198e+01                   4
C14H9                   C  14H   9          G    298.15   3500.00 1380.00      1
 2.51054802e+01 4.12375730e-02-1.71094078e-05 3.35330064e-09-2.55891906e-13    2
 4.20489545e+04-1.12231128e+02-1.15966331e+01 1.47620510e-01-1.32743035e-04    3
 5.92149564e-08-1.03757571e-11 5.21787378e+04 7.66564976e+01                   4
C16H10                  C  16H  10          G    200.00   3500.00 1560.00      1
 3.81807346e+01 2.83119223e-02-6.73305412e-06 1.57165249e-10 8.21178664e-14    2
 9.09208909e+03-1.88517714e+02-1.17161985e+01 1.56252776e-01-1.29753106e-04    3
 5.27298370e-08-8.34298979e-12 2.46599322e+04 7.43946040e+01                   4
C16H9                   C  16H   9          G    300.00   3500.00 1240.00      1
 1.61933978e+01 6.96117135e-02-3.71054120e-05 9.43826012e-09-9.32515878e-13    2
 4.61008358e+04-6.54256239e+01-1.33382684e+01 1.64875153e-01-1.52343444e-04    3
 7.13941910e-08-1.34236310e-11 5.34246890e+04 8.34001921e+01                   4
C6H5C2H4C6H5            C  14H  14          G    300.00   3500.00 1170.00      1
 6.79293353e+00 9.36089894e-02-5.25184355e-05 1.38852184e-08-1.40951794e-12    2
 1.04787082e+04-8.65156283e+00-1.16088786e+01 1.56521168e-01-1.33175074e-04    3
 5.98434171e-08-1.12296459e-11 1.47847322e+04 8.30156968e+01                   4
C18H10                  C  18H  10          G    300.00   3500.00 1430.00      1
 3.55205899e+01 2.97059393e-02-5.18578691e-06-7.74972602e-10 2.05763862e-13    2
 1.13998056e+04-1.72584615e+02-1.43149505e+01 1.69106052e-01-1.51409682e-04    3
 6.73946752e-08-1.17120067e-11 2.56527701e+04 8.56679583e+01                   4
C18H9                   C  18H   9          G    300.00   3500.00 1110.00      1
 1.00826780e+01 9.26185738e-02-5.34378516e-05 1.44603235e-08-1.49786389e-12    2
 4.90427510e+04-3.41228885e+01-1.54340436e+01 1.84570724e-01-1.77697514e-04    3
 8.90907512e-08-1.83065188e-11 5.47074632e+04 9.16434687e+01                   4
LC6H5                   C   6H   5          G    300.00   3500.00 1140.00      1
 1.23076076e+01 1.68261951e-02-6.51181367e-06 1.21158890e-09-8.99428205e-14    2
 5.89425072e+04-3.55373249e+01 1.67614161e-01 5.94226633e-02-6.25597981e-05    3
 3.39881880e-08-7.27779349e-12 6.17104257e+04 2.46218080e+01                   4
C6H2                    C   6H   2          G    200.00   3500.00  700.00      1
 9.95239961e+00 1.43744770e-02-7.32585546e-06 1.80931772e-09-1.74471745e-13    2
 8.06473020e+04-2.49945457e+01-5.39476453e-01 7.43280545e-02-1.35797807e-04    3
 1.24163557e-07-4.38724145e-11 8.21161647e+04 2.18805021e+01                   4
C6H3                    C   6H   3          G    300.00   3500.00 1320.00      1
 1.19194523e+01 1.16137832e-02-4.19264521e-06 6.84693068e-10-4.17887563e-14    2
 8.26280760e+04-3.29876543e+01 4.46601449e+00 3.41999583e-02-2.98587533e-05    3
 1.36473739e-08-2.49684195e-12 8.45957836e+04 5.04018538e+00                   4
C6H4                    C   6H   4          G    300.00   3500.00 1360.00      1
 1.74447675e+01 6.21306704e-03-9.80963831e-07 8.00594547e-11-2.88320672e-15    2
 5.49568894e+04-6.59208083e+01-1.17305610e+00 6.09713718e-02-6.13761529e-05    3
 2.96855443e-08-5.44506792e-12 6.00209374e+04 2.96241244e+01                   4
C8H2                    C   8H   2          G    300.00   3500.00 1060.00      1
 1.62719352e+01 9.99874483e-03-2.93037073e-06 2.89537319e-10 2.52408504e-16    2
 1.07885460e+05-5.89733616e+01 1.87361690e-01 7.06952486e-02-8.88216497e-05    3
 5.43092096e-08-1.27402363e-11 1.11295389e+05 1.95626384e+01                   4
C18H14                  H  14C  18          G    100.00   3500.00  700.00      1
-8.78909816e+00 1.54177573e-01-9.84392858e-05 2.89551422e-08-3.12416385e-12    2
 3.49494076e+04 6.52592557e+01-7.00582263e+00 1.43987427e-01-7.66032589e-05    3
 8.15892605e-09 4.30305619e-12 3.46997490e+04 5.72920318e+01                   4
BIN1A                   C  20H  16          G    300.00   3500.00 1410.00      1
 4.18189976e+01 5.54173538e-02-1.89314485e-05 2.76164872e-09-1.34640910e-13    2
-3.16800426e+03-2.10125738e+02-1.45702439e+01 2.15386833e-01-1.89111746e-04    3
 8.32251462e-08-1.44012185e-11 1.27337618e+04 8.12945187e+01                   4
BIN1B                   C  20H  10          G    300.00   3500.00 1430.00      1
 3.76362494e+01 4.45434540e-02-1.43416602e-05 1.85353053e-09-6.45805559e-14    2
-9.82259725e+02-1.87789164e+02-1.59101514e+01 1.94323596e-01-1.71453697e-04    3
 7.50992355e-08-1.28697737e-11 1.43320109e+04 8.96934466e+01                   4
FC10H10                 C  10H  10          G    300.00   3500.00 1800.00      1
 1.82592698e+01 4.15934215e-02-1.83631831e-05 3.88491134e-09-3.27420807e-13    2
 4.39687820e+03-8.23923220e+01-1.14588964e+01 1.07633791e-01-7.33968243e-05    3
 2.42677414e-08-3.15836943e-12 1.50954180e+04 7.84485932e+01                   4
C6H5C2H4                C   8H   9          G    200.00   3500.00 1530.00      1
 1.90733241e+01 2.32393227e-02-7.04814668e-06 8.06136144e-10-1.68209988e-14    2
 1.95612163e+04-7.66267161e+01-3.58296948e+00 8.24714629e-02-6.51188723e-05    3
 2.61092846e-08-4.15132238e-12 2.64940422e+04 4.23117947e+01                   4
RMCYC6                  C   7H  13          G    300.00   3500.00 1800.00      1
 1.73339062e+01 3.85260822e-02-1.58310821e-05 3.15191459e-09-2.53163787e-13    2
-5.89957979e+03-7.33836419e+01-9.95790328e+00 9.91745477e-02-6.63714701e-05    3
 2.18705768e-08-2.85297798e-12 3.92547162e+03 7.43253244e+01                   4
MCYC6                   C   7H  14          G    300.00   3500.00 1800.00      1
 1.67194568e+01 4.36180644e-02-1.87773363e-05 3.92059022e-09-3.26702984e-13    2
-2.91866300e+04-7.40611877e+01-1.01006358e+01 1.03218270e-01-6.84441744e-05    3
 2.23157154e-08-2.88158149e-12-1.95313967e+04 7.10947481e+01                   4
TMBENZ                  C   9H  12          G    300.00   3500.00 1800.00      1
 1.47576861e+01 4.50315825e-02-1.97554195e-05 4.21197817e-09-3.57314917e-13    2
-1.09025839e+04-5.35378398e+01-2.75522789e+00 8.39491691e-02-5.21867417e-05    3
 1.62235790e-08-2.02559281e-12-4.59793488e+03 4.12457040e+01                   4
NPBENZ                  C   9H  12          G    300.00   3500.00 1600.00      1
 1.88963371e+01 3.80090295e-02-1.52789389e-05 2.95630099e-09-2.27699217e-13    2
-8.96605283e+03-7.62711275e+01-5.58650157e+00 9.92161261e-02-7.26605920e-05    3
 2.68653231e-08-3.96348393e-12-1.13154446e+03 5.33514397e+01                   4
RC9H11                  C   9H  11          G    300.00   3500.00 1800.00      1
 1.94777671e+01 3.52558916e-02-1.42493230e-05 2.76058348e-09-2.13045169e-13    2
 6.10938819e+03-7.94713741e+01-1.83523003e+00 8.26181075e-02-5.37178363e-05    3
 1.73785513e-08-2.24331848e-12 1.37820672e+04 3.58790126e+01                   4
DIBZFUR                 C  12H   8O   1     G    300.00   3500.00 1410.00      1
 2.49525256e+01 3.24730728e-02-1.15459374e-05 1.79679053e-09-9.97833648e-14    2
-5.30753652e+03-1.13355893e+02-1.16970901e+01 1.36443614e-01-1.22152896e-04    3
 5.40932248e-08-9.37220079e-12 5.02765510e+03 7.60497478e+01                   4
BZFUR                   C   8H   6O   1     G    300.00   3500.00 1380.00      1
 1.64578334e+01 2.37623566e-02-8.52218596e-06 1.36123709e-09-7.97159879e-14    2
-5.90596973e+03-6.59480382e+01-8.70136948e+00 9.66875824e-02-8.77887357e-05    3
 3.96542563e-08-7.01685715e-12 1.03797027e+03 6.35339364e+01                   4
ODECAL                  C  10H  18          G    300.00   3500.00 1800.00      1
 2.82109941e+01 4.74108396e-02-1.82963852e-05 3.42084161e-09-2.57817125e-13    2
-2.68355230e+04-1.31410203e+02-1.02710769e+01 1.32926553e-01-8.95594797e-05    3
 2.98145803e-08-3.92361417e-12-1.29819774e+04 7.68627930e+01                   4
DECALIN                 C  10H  18          G    300.00   3500.00 1750.00      1
 2.70110296e+01 4.68748171e-02-1.63895490e-05 2.62563687e-09-1.59789734e-13    2
-3.79226289e+04-1.35167747e+02-1.45870783e+01 1.41956207e-01-9.78878828e-05    3
 3.36726212e-08-4.59507321e-12-2.33632912e+04 8.87980358e+01                   4
TETRALIN                C  10H  12          G    300.00   3500.00 1650.00      1
 2.40250678e+01 3.45031690e-02-1.26565536e-05 2.20632463e-09-1.51941206e-13    2
-9.85314330e+03-1.11161769e+02-1.00807336e+01 1.17183900e-01-8.78208542e-05    3
 3.25757390e-08-4.75336763e-12 1.40177116e+03 7.04583499e+01                   4
DCYC5                   C  10H  16          G    300.00   3500.00 1750.00      1
 2.70110296e+01 4.68748172e-02-1.63895490e-05 2.62563687e-09-1.59789734e-13    2
-3.79226289e+04-1.35167747e+02-1.45870783e+01 1.41956207e-01-9.78878828e-05    3
 3.36726212e-08-4.59507321e-12-2.33632912e+04 8.87980358e+01                   4
RTETRALIN               C  10H  11          G    300.00   3500.00 1800.00      1
 2.92428061e+01 2.67835938e-02-9.17249483e-06 1.42952537e-09-8.46466190e-14    2
 3.95646505e+03-1.44540610e+02-1.09331574e+01 1.16063513e-01-8.35724273e-05    3
 2.89850559e-08-3.91180364e-12 1.84198119e+04 7.29000859e+01                   4
RTETRAOO                C  10H  11O   2     G    300.00   3500.00 1800.00      1
 5.34619031e+01-7.89283130e-03 1.09697206e-05-3.89489829e-09 4.38586293e-13    2
-1.76924159e+04-2.71823424e+02-1.36343924e+01 1.41210048e-01-1.13282678e-04    3
 4.21245088e-08-5.95299802e-12 6.46225047e+03 9.13157248e+01                   4
RDECALIN                C  10H  17          G    300.00   3500.00 1800.00      1
 2.85620333e+01 4.11366392e-02-1.36024110e-05 2.01592783e-09-1.09376626e-13    2
-1.53025063e+04-1.39641687e+02-1.39601308e+01 1.35630337e-01-9.23471594e-05    3
 3.11806495e-08-4.16003241e-12 5.47278060e+00 9.04971362e+01                   4
RODECA                  C  10H  17          G    300.00   3500.00 1800.00      1
 2.85620333e+01 4.11366392e-02-1.36024110e-05 2.01592783e-09-1.09376626e-13    2
-1.53025063e+04-1.39641687e+02-1.39601308e+01 1.35630337e-01-9.23471594e-05    3
 3.11806495e-08-4.16003241e-12 5.47278060e+00 9.04971362e+01                   4
NC10H22                 C  10H  22          G    300.00   3500.00 1800.00      1
 2.92878918e+01 5.29920990e-02-1.98404553e-05 3.55616370e-09-2.54281184e-13    2
-4.56232379e+04-1.22752047e+02-2.17870143e+00 1.22917862e-01-7.81119243e-05    3
 2.51381892e-08-3.25178473e-12-3.42952643e+04 4.75517200e+01                   4
NC10H21                 C  10H  21          G    300.00   3500.00 1800.00      1
 2.63212692e+01 5.52219738e-02-2.21266526e-05 4.33498891e-09-3.42316503e-13    2
-2.10175171e+04-1.03192977e+02-1.81057271e+00 1.17737178e-01-7.42226562e-05    3
 2.36298050e-08-3.02215208e-12-1.08900540e+04 4.90624204e+01                   4
C10H10                  C  10H  10          G    300.00   3500.00 1800.00      1
 1.82592698e+01 4.15934215e-02-1.83631831e-05 3.88491134e-09-3.27420807e-13    2
 4.39687820e+03-8.23923220e+01-1.14588964e+01 1.07633791e-01-7.33968243e-05    3
 2.42677414e-08-3.15836943e-12 1.50954180e+04 7.84485932e+01                   4
NC12H25                 C  12H  25          G    300.00   3500.00 1800.00      1
 3.17005579e+01 6.61544325e-02-2.66295230e-05 5.21804510e-09-4.10998519e-13    2
-2.88525898e+04-1.31607624e+02-2.06085145e+00 1.41179787e-01-8.91506513e-05    3
 2.83740186e-08-3.62710594e-12-1.66984825e+04 5.11161660e+01                   4
IC16H33                 C  16H  33          G    300.00   3500.00 1650.00      1
 5.11453588e+01 7.53296743e-02-2.79263242e-05 4.92908201e-09-3.44364401e-13    2
-5.61938874e+04-2.43048234e+02-8.95216176e+00 2.21020633e-01-1.60372651e-04    3
 5.84427492e-08-8.45249580e-12-3.63617056e+04 7.69829165e+01                   4
NC16H33                 C  16H  33          G    300.00   3500.00 1800.00      1
 4.66278371e+01 8.00212238e-02-3.03236334e-05 5.55903617e-09-4.09822554e-13    2
-4.61545210e+04-2.04019480e+02-3.22413374e+00 1.90803381e-01-1.22642098e-04    3
 3.97510601e-08-5.15871477e-12-2.82078115e+04 6.57897857e+01                   4
NC10H19                 C  10H  19          G    300.00   3500.00 1800.00      1
 9.88287390e+00 2.86275350e-02-1.23662428e-05 2.58308509e-09-2.14520963e-13    2
 7.14211639e+03-2.81379758e+01-9.61360662e-01 5.27258341e-02-3.24481586e-05    3
 1.00208317e-08-1.24754133e-12 1.10460408e+04 3.05532839e+01                   4
NC12H26                 C  12H  26          G    300.00   3500.00 1800.00      1
 3.61414094e+01 6.11045883e-02-2.24641073e-05 3.93182441e-09-2.73349363e-13    2
-5.40359186e+04-1.56831960e+02-2.66627705e+00 1.47343892e-01-9.43301934e-05    3
 3.05488933e-08-3.97016449e-12-4.00651514e+04 5.32033350e+01                   4
IC16H34                 C  16H  34          G    300.00   3500.00 1590.00      1
 4.72524599e+01 8.54680758e-02-3.36612723e-05 6.38202030e-09-4.82094888e-13    2
-7.78744142e+04-2.24182950e+02-9.93612249e+00 2.29338723e-01-1.69388298e-04    3
 6.32906266e-08-9.42998896e-12-5.96884450e+04 7.82391931e+01                   4
NC16H34                 C  16H  34          G    300.00   3500.00 1800.00      1
 4.98210237e+01 7.73881688e-02-2.77557896e-05 4.69678103e-09-3.12959243e-13    2
-7.08514663e+04-2.24842855e+02-3.64057977e+00 1.96191732e-01-1.26758759e-04    3
 4.13645475e-08-5.40570458e-12-5.16052891e+04 6.45024954e+01                   4
NC10H20                 C  10H  20          G    300.00   3500.00 1800.00      1
 2.82971791e+01 4.89478938e-02-1.82737062e-05 3.23575201e-09-2.26811842e-13    2
-3.12534582e+04-1.16784058e+02-2.31417710e+00 1.16973130e-01-7.49614029e-05    3
 2.42311952e-08-3.14284563e-12-2.02333700e+04 4.88909878e+01                   4
IC12H26                 C  12H  26          G    300.00   3500.00 1800.00      1
 3.61414094e+01 6.11045883e-02-2.24641073e-05 3.93182441e-09-2.73349363e-13    2
-5.40359186e+04-1.56831960e+02-2.66627705e+00 1.47343892e-01-9.43301934e-05    3
 3.05488933e-08-3.97016449e-12-4.00651514e+04 5.32033350e+01                   4
IC12H25                 C  12H  25          G    300.00   3500.00 1800.00      1
 3.17005579e+01 6.61544325e-02-2.66295230e-05 5.21804510e-09-4.10998519e-13    2
-2.88525898e+04-1.31607624e+02-2.06085145e+00 1.41179787e-01-8.91506513e-05    3
 2.83740186e-08-3.62710594e-12-1.66984825e+04 5.11161660e+01                   4
C10H16                  C  10H  16          G    300.00   3500.00 1800.00      1
 2.89286921e+01 4.33698641e-02-1.66040771e-05 3.00058011e-09-2.14826944e-13    2
-2.62354027e+04-1.44986840e+02-1.64117649e+01 1.44126435e-01-1.00567886e-04    3
 3.40982872e-08-4.53395293e-12-9.91283823e+03 1.00405171e+02                   4
C10H15                  C  10H  15          G    300.00   3500.00 1770.00      1
 3.20501672e+01 3.53882361e-02-1.22004701e-05 1.87186214e-09-1.05121248e-13    2
-9.38259390e+03-1.63611897e+02-1.67888481e+01 1.45758892e-01-1.05734924e-04    3
 3.71014118e-08-5.08104634e-12 7.90641753e+03 9.98941988e+01                   4
C6H5C4H9                C  10H  14          G    300.00   3500.00 1620.00      1
 2.20508088e+01 4.25105888e-02-1.68597965e-05 3.21476378e-09-2.44036713e-13    2
-1.30455855e+04-9.17623601e+01-5.81141602e+00 1.11306205e-01-8.05594416e-05    3
 2.94286095e-08-4.28938328e-12-4.01822468e+03 5.60982344e+01                   4
RC6H5C4H8               C  10H  13          G    300.00   3500.00 1650.00      1
 2.28150862e+01 3.94891782e-02-1.56943357e-05 2.97948809e-09-2.24328827e-13    2
 4.22313026e+03-9.69374623e+01-3.49464028e+00 1.03270333e-01-7.36772040e-05    3
 2.64069096e-08-3.77393815e-12 1.29053400e+04 4.31670204e+01                   4
C6H5C4H7-3              C  10H  12          G    300.00   3500.00 1480.00      1
 1.62604546e+01 4.74926138e-02-2.11208270e-05 4.52915802e-09-3.83727993e-13    2
 2.53220324e+03-5.97390118e+01-5.26848595e+00 1.05678940e-01-8.00934545e-05    3
 3.10934047e-08-4.87093182e-12 8.90476965e+03 5.25659324e+01                   4
CH2OHCH2OH              C   2H   6O   2     G    300.00   3500.00 1510.00      1
 8.58229286e+00 1.47365725e-02-4.87454255e-06 7.03407966e-10-3.54291380e-14    2
-5.09140292e+04-1.61663169e+01-4.19778978e-01 3.85831204e-02-2.85631663e-05    3
 1.11619615e-08-1.76697774e-12-4.81954035e+04 3.09733167e+01                   4
GLYCEROL                C   3H   8O   3     G    300.00   3500.00 1260.00      1
 1.38765805e+01 2.06689859e-02-7.56631173e-06 1.26540495e-09-8.07916650e-14    2
-7.51651919e+04-3.83652419e+01 3.56065369e+00 5.34179600e-02-4.65531857e-05    3
 2.18933806e-08-4.17364397e-12-7.25655783e+04 1.37872736e+01                   4
C3H4O3                  C   3H   4O   3     G    300.00   3500.00 1710.00      1
 1.37242810e+01 1.08811110e-02-3.70124855e-06 5.78901441e-10-3.43205819e-14    2
-5.77802807e+04-3.99570073e+01 2.17563103e+00 3.78954970e-02-2.73980784e-05    3
 9.81743158e-09-1.38498288e-12-5.38306424e+04 2.19543274e+01                   4
FURFURAL                C   5H   4O   2     G    300.00   3500.00 1430.00      1
 1.05158963e+01 2.23224229e-02-1.09267096e-05 2.56683236e-09-2.34844996e-13    2
-2.33303219e+04-2.94000375e+01-1.81996645e+00 5.68283326e-02-4.71217198e-05    3
 1.94409630e-08-3.18486783e-12-1.98022652e+04 3.45255921e+01                   4
FURAN                   C   4H   4O   1     G    300.00   3500.00 1250.00      1
 8.37486468e+00 1.95634451e-02-9.90167118e-06 2.37694381e-09-2.20517697e-13    2
-9.41817580e+03-2.52053385e+01-7.59507782e+00 7.06672611e-02-7.12262504e-05    3
 3.50833860e-08-6.76180614e-12-5.42569018e+03 5.54039923e+01                   4
CH2CCHCHO               C   4H   4O   1     G    300.00   3500.00 1590.00      1
 1.05858550e+01 1.29956017e-02-4.76361254e-06 7.49449812e-10-3.96847799e-14    2
 3.10513348e+03-2.93262371e+01 1.05972039e+00 3.69607201e-02-2.73722149e-05    3
 1.02289476e-08-1.53017186e-12 6.13444428e+03 2.10494483e+01                   4
C4H3O                   C   4H   3O   1     G    300.00   3500.00 1240.00      1
 8.44125907e+00 1.62911135e-02-8.34126433e-06 2.01436765e-09-1.87394602e-13    2
 1.94535776e+04-2.27855079e+01-5.90872254e+00 6.25813768e-02-6.43375505e-05    3
 3.21198979e-08-6.25705795e-12 2.30123730e+04 4.95317027e+01                   4
MEFU2                   C   5H   6O   1     G    300.00   3500.00 1260.00      1
 5.16398170e+00 3.29529080e-02-1.68209195e-05 4.03716052e-09-3.55511368e-13    2
-1.31841670e+04-2.67616715e+00-3.74149805e+00 6.12242723e-02-5.04773056e-05    3
 2.18447722e-08-3.88876765e-12-1.09399861e+04 4.23457855e+01                   4
DMF                     C   6H   8O   1     G    300.00   3500.00 1590.00      1
 1.38889506e+01 2.49736923e-02-8.98421019e-06 1.42738237e-09-7.97717940e-14    2
-2.20872034e+04-4.94041110e+01-2.31533181e+00 6.57391826e-02-4.74422199e-05    3
 1.75523340e-08-2.61514155e-12-1.69342416e+04 3.62866615e+01                   4
DMF-3YL                 C   6H   7O   1     G    300.00   3500.00 1620.00      1
 1.41703395e+01 2.18230092e-02-7.69511406e-06 1.17891300e-09-6.12376633e-14    2
 1.19557792e+04-4.86583490e+01-1.12307985e+00 5.95845385e-02-4.26594930e-05    3
 1.55675463e-08-2.28170577e-12 1.69108471e+04 3.25015044e+01                   4
C6H10O5                 C   6H  10O   5     G    300.00   3500.00 1220.00      1
 1.54889719e+01 4.96354386e-02-2.45944508e-05 5.82332583e-09-5.35665861e-13    2
-1.09180509e+05-4.81819838e+01-7.95116462e+00 1.26488345e-01-1.19085729e-04    3
 5.74579043e-08-1.11165221e-11-1.03461116e+05 6.95642163e+01                   4
C6H8O4                  C   6H   8O   4     G    300.00   3500.00 1300.00      1
 1.58073709e+01 3.77998882e-02-1.77241312e-05 3.97560136e-09-3.49009860e-13    2
-7.78788467e+04-5.15128322e+01-4.55493836e+00 1.00453147e-01-9.00163533e-05    3
 4.10485358e-08-7.47842033e-12-7.25846463e+04 5.20658817e+01                   4
C6H6O3                  C   6H   6O   3     G    300.00   3500.00 1770.00      1
 1.98638073e+01 1.79335016e-02-5.95408858e-06 8.93593938e-10-4.95459879e-14    2
-4.95264845e+04-7.44496694e+01 7.10718581e-01 6.12173180e-02-4.26352889e-05    3
 1.47094886e-08-2.00094354e-12-4.27462910e+04 2.88889342e+01                   4
C5H8O4                  C   5H   8O   4     G    300.00   3500.00 1230.00      1
 1.19601536e+01 3.99450842e-02-1.95947372e-05 4.60940116e-09-4.22302288e-13    2
-8.26385858e+04-2.91875209e+01-6.95683232e+00 1.01463738e-01-9.46174852e-05    3
 4.52721372e-08-8.68708604e-12-7.79850073e+04 6.59920851e+01                   4
CATECHOL                C   6H   6O   2     G    300.00   3500.00 1150.00      1
 1.43499798e+01 2.44086034e-02-1.04210955e-05 2.01938915e-09-1.47232753e-13    2
-3.94515399e+04-4.76262861e+01-5.49815264e+00 9.34455857e-02-1.00469333e-04    3
 5.42212661e-08-1.14954669e-11-3.48864694e+04 5.09034930e+01                   4
GUAIACOL                C   7H   8O   2     G    300.00   3500.00 1000.00      1
 9.99301702e+00 4.50609511e-02-2.36180854e-05 5.74986028e-09-5.33615163e-13    2
-3.55531885e+04-2.30989094e+01-7.52910625e+00 1.15149444e-01-1.28750825e-04    3
 7.58383534e-08-1.80557384e-11-3.20487639e+04 6.14352066e+01                   4
SALICALD                C   7H   6O   2     G    300.00   3500.00 1580.00      1
 2.23242869e+01 1.54051239e-02-2.83991520e-06-4.41655604e-10 1.22876781e-13    2
-3.64536802e+04-8.95534660e+01-5.00623399e+00 8.45963160e-02-6.85277558e-05    3
 2.72747329e-08-4.26262772e-12-2.78172356e+04 5.48021581e+01                   4
VANILLIN                C   8H   8O   3     G    300.00   3500.00 1260.00      1
 1.36544657e+01 4.84143206e-02-2.42641773e-05 5.50487741e-09-4.76001842e-13    2
-5.18855417e+04-3.54575763e+01-4.86637434e+00 1.07210638e-01-9.42597934e-05    3
 4.25395949e-08-7.82416008e-12-4.72182901e+04 5.81751540e+01                   4
C8H6O3                  C   8H   6O   3     G    300.00   3500.00 1000.00      1
 4.59308938e+00 6.23299053e-02-3.47374653e-05 8.74937512e-09-8.39789340e-13    2
-4.48191760e+04 1.51136268e+01-8.47052157e+00 1.14584349e-01-1.13119131e-04    3
 6.10038189e-08-1.39034003e-11-4.22064538e+04 7.81379982e+01                   4
C6H5OCH3                C   7H   8O   1     G    300.00   3500.00 1380.00      1
 1.25085136e+01 3.49906122e-02-1.63096082e-05 3.64836833e-09-3.19988393e-13    2
-1.52038795e+04-4.20406498e+01-5.29461551e+00 8.65938851e-02-7.24001222e-05    3
 3.07452350e-08-5.22884105e-12-1.02902159e+04 4.95832512e+01                   4
C7H6O3                  C   7H   6O   3     G    300.00   3500.00 1000.00      1
 9.61003482e+00 4.63126508e-02-2.49854466e-05 6.23131070e-09-5.96782041e-13    2
-5.28813088e+04-1.46625767e+01-7.07010661e+00 1.13033217e-01-1.25066295e-04    3
 7.29518764e-08-1.72769235e-11-4.95452805e+04 6.58094637e+01                   4
RC7H5O3                 C   7H   5O   3     G    300.00   3500.00 1000.00      1
 1.03519979e+01 4.06949751e-02-2.16398121e-05 5.16863286e-09-4.69580368e-13    2
-3.48541025e+04-1.78724723e+01-6.94106369e+00 1.09867221e-01-1.25398181e-04    3
 7.43408790e-08-1.77626419e-11-3.13954902e+04 6.55565533e+01                   4
C24H28O4                C  24H  28O   4     G    300.00   3500.00 1080.00      1
 1.29252083e+01 8.11297204e-02-4.64957343e-05 1.23575596e-08-1.22239418e-12    2
-7.66058401e+03-2.94388917e+00 3.08710551e+00 1.17567138e-01-9.71032588e-05    3
 4.35967723e-08-8.45369342e-12-5.53555381e+03 4.52764204e+01                   4
C6H4O                   C   6H   4O   1     G    300.00   3500.00 1320.00      1
 1.34428169e+01 1.79658729e-02-6.67332776e-06 1.12237516e-09-7.10809492e-14    2
 1.54076839e+04-4.72500521e+01-4.80707079e+00 7.32685627e-02-6.95172935e-05    3
 3.28617518e-08-6.08232653e-12 2.02256542e+04 4.58618545e+01                   4
RSALICPH                C   7H   5O   2     G    300.00   3500.00 1000.00      1
 6.00653618e+00 4.55336023e-02-2.51852438e-05 6.39158463e-09-6.19568356e-13    2
 4.68000597e+02 2.82366668e+00-8.00629363e+00 1.01584922e-01-1.09262223e-04    3
 6.24429039e-08-1.46323982e-11 3.27056656e+03 7.04274704e+01                   4
RGUAIPH                 C   7H   7O   2     G    300.00   3500.00 1000.00      1
 1.03288605e+01 4.15815436e-02-2.20221230e-05 5.39151185e-09-5.01575209e-13    2
-4.91455279e+03-2.20047760e+01-7.23884832e+00 1.11852379e-01-1.27428376e-04    3
 7.56623473e-08-1.80692841e-11-1.40101102e+03 6.27492641e+01                   4
RANISPH                 C   7H   7O   1     G    300.00   3500.00 1000.00      1
 6.14038338e+00 4.52741698e-02-2.46495239e-05 6.30633007e-09-6.15603035e-13    2
 1.78813933e+04-4.35386646e+00-8.02841875e+00 1.01949378e-01-1.09662337e-04    3
 6.29815386e-08-1.47844052e-11 2.07151538e+04 6.40024135e+01                   4
RCATEPH                 C   6H   5O   2     G    300.00   3500.00 1000.00      1
 1.18218909e+01 2.70911128e-02-1.34162451e-05 3.08575096e-09-2.72412002e-13    2
-7.82412457e+03-3.10506064e+01-7.41421160e+00 1.04035523e-01-1.28832860e-04    3
 8.00301608e-08-1.95085145e-11-3.97690408e+03 6.17524685e+01                   4
BIN1C                   C  20H   5          G    300.00   3500.00 1390.00      1
 3.44720380e+01 3.60523047e-02-1.05663116e-05 1.05180871e-09 2.58274737e-15    2
-8.53118933e+03-1.83953590e+02-1.67831316e+01 1.83549196e-01-1.69735618e-04    3
 7.73920039e-08-1.37276682e-11 5.71774783e+03 8.02014943e+01                   4
BIN2A                   C  40H  31          G    300.00   3500.00 1380.00      1
 8.09167423e+01 1.12943669e-01-3.95771786e-05 6.05002182e-09-3.25324880e-13    2
-1.79932662e+03-4.04172972e+02-3.17321030e+01 4.39462062e-01-3.94488475e-04    3
 1.77504754e-07-3.13859648e-11 2.92917547e+04 1.75574924e+02                   4
BIN2B                   C  40H  16          G    300.00   3500.00 1410.00      1
 7.17877214e+01 8.40138218e-02-2.68733543e-05 3.42345855e-09-1.13355144e-13    2
-8.39424360e+03-3.65933272e+02-3.29263051e+01 3.81074890e-01-3.42895767e-04    3
 1.52843039e-07-2.66061886e-11 2.11351119e+04 1.75230037e+02                   4
BIN2C                   C  40H   8          G    300.00   3500.00 1390.00      1
 6.81202262e+01 6.75222092e-02-1.89112417e-05 1.59405249e-09 5.05762487e-14    2
-2.22065321e+04-3.64909286e+02-3.46582201e+01 3.63287522e-01-3.38082443e-04    3
 1.54673765e-07-2.74817462e-11 6.36587595e+03 1.64782634e+02                   4
BIN3A                   C  80H  60          G    300.00   3500.00 1360.00      1
 1.60725588e+02 2.23424535e-01-7.78333867e-05 1.17513969e-08-6.14855228e-13    2
-1.27263143e+03-8.20183331e+02-6.32696159e+01 8.82233959e-01-8.04461428e-04    3
 3.67941613e-07-6.60909979e-11 5.96540641e+04 3.29339146e+02                   4
BIN3B                   C  80H  24          G    300.00   3500.00 1400.00      1
 1.39875812e+02 1.51591568e-01-4.58194656e-05 5.02696436e-09-6.37152147e-14    2
-3.05860818e+04-7.30660869e+02-6.75753698e+01 7.44309230e-01-6.80874104e-04    3
 3.07433935e-07-5.40649600e-11 2.75002491e+04 3.39972729e+02                   4
BIN3C                   C  80H   8          G    300.00   3500.00 1380.00      1
 1.32666452e+02 1.18391629e-01-2.97594453e-05 1.33141073e-09 2.67779755e-13    2
-5.82681507e+04-7.29323376e+02-7.10761933e+01 7.08950020e-01-6.71670740e-04    3
 3.11433486e-07-5.59101324e-11-2.03518064e+03 3.19239256e+02                   4
BIN1AJ                  C  20H  15          G    300.00   3500.00 1410.00      1
 4.18189976e+01 5.54173538e-02-1.89314485e-05 2.76164872e-09-1.34640910e-13    2
 5.68319957e+04-2.10125738e+02-1.45702439e+01 2.15386833e-01-1.89111746e-04    3
 8.32251462e-08-1.44012185e-11 7.27337618e+04 8.12945187e+01                   4
BIN1BJ                  C  20H   9          G    300.00   3500.00 1430.00      1
 3.76362494e+01 4.45434540e-02-1.43416602e-05 1.85353053e-09-6.45805559e-14    2
 5.90177403e+04-1.87789164e+02-1.59101514e+01 1.94323596e-01-1.71453697e-04    3
 7.50992355e-08-1.28697737e-11 7.43320109e+04 8.96934466e+01                   4
BIN1CJ                  C  20H   4          G    300.00   3500.00 1390.00      1
 3.44720380e+01 3.60523047e-02-1.05663116e-05 1.05180871e-09 2.58274737e-15    2
 5.14688106e+04-1.83953590e+02-1.67831316e+01 1.83549196e-01-1.69735618e-04    3
 7.73920039e-08-1.37276682e-11 6.57177478e+04 8.02014943e+01                   4
BIN2AJ                  C  40H  30          G    300.00   3500.00 1380.00      1
 8.09167423e+01 1.12943669e-01-3.95771786e-05 6.05002182e-09-3.25324880e-13    2
 5.82006734e+04-4.04172972e+02-3.17321030e+01 4.39462062e-01-3.94488475e-04    3
 1.77504754e-07-3.13859648e-11 8.92917547e+04 1.75574924e+02                   4
BIN2BJ                  C  40H  15          G    300.00   3500.00 1410.00      1
 7.17877214e+01 8.40138218e-02-2.68733543e-05 3.42345855e-09-1.13355144e-13    2
 5.16057564e+04-3.65933272e+02-3.29263051e+01 3.81074890e-01-3.42895767e-04    3
 1.52843039e-07-2.66061886e-11 8.11351119e+04 1.75230037e+02                   4
BIN2CJ                  C  40H   7          G    300.00   3500.00 1390.00      1
 6.81202262e+01 6.75222092e-02-1.89112417e-05 1.59405249e-09 5.05762487e-14    2
 3.77934679e+04-3.64909286e+02-3.46582201e+01 3.63287522e-01-3.38082443e-04    3
 1.54673765e-07-2.74817462e-11 6.63658759e+04 1.64782634e+02                   4
BIN3AJ                  C  80H  59          G    300.00   3500.00 1360.00      1
 1.60725588e+02 2.23424535e-01-7.78333867e-05 1.17513969e-08-6.14855228e-13    2
 5.87273686e+04-8.20183331e+02-6.32696159e+01 8.82233959e-01-8.04461428e-04    3
 3.67941613e-07-6.60909979e-11 1.19654064e+05 3.29339146e+02                   4
BIN3BJ                  C  80H  23          G    300.00   3500.00 1400.00      1
 1.39875812e+02 1.51591568e-01-4.58194656e-05 5.02696436e-09-6.37152147e-14    2
 2.94139182e+04-7.30660869e+02-6.75753698e+01 7.44309230e-01-6.80874104e-04    3
 3.07433935e-07-5.40649600e-11 8.75002491e+04 3.39972729e+02                   4
BIN3CJ                  C  80H   7          G    300.00   3500.00 1380.00      1
 1.32666452e+02 1.18391629e-01-2.97594453e-05 1.33141073e-09 2.67779755e-13    2
 1.73184933e+03-7.29323376e+02-7.10761933e+01 7.08950020e-01-6.71670740e-04    3
 3.11433486e-07-5.59101324e-11 5.79648194e+04 3.19239256e+02                   4
BIN4AJ                                      G    300.00   3500.00 1330.00      1&
C 160.00 H 115.00 
 3.13388326e+02 4.53632950e-01-1.61287498e-04 2.52639660e-08-1.42054928e-12    2
 6.43001833e+04-1.63197350e+03-1.27820190e+02 1.78057585e+00-1.65783965e-03    3
 7.75415418e-07-1.42426461e-10 1.81661648e+05 6.22425921e+02                   4
BIN4BJ                                      G    300.00   3500.00 1390.00      1&
C 160.00 H 31.00 
 2.72480905e+02 2.70088841e-01-7.56449720e-05 6.37621196e-09 2.02304741e-13    2
-2.88261298e+04-1.45963715e+03-1.38632883e+02 1.45315010e+00-1.35232978e-03    3
 6.18695067e-07-1.09926986e-10 8.54635032e+04 6.59130542e+02                   4
BIN4CJ                                      G    300.00   3500.00 1370.00      1&
C 160.00 H 9.00 
 2.59057611e+02 2.31346303e-01-5.83745085e-05 2.71298902e-09 5.07830703e-13    2
-6.54530912e+04-1.43847454e+03-1.44192320e+02 1.40871836e+00-1.34746801e-03    3
 6.30009095e-07-1.13962262e-10 4.50373899e+04 6.33920690e+02                   4
BIN5AJ                                      G    300.00   3500.00 1310.00      1&
C 320.00 H 223.00 
 6.22157978e+02 8.96699580e-01-3.17277804e-04 4.92175274e-08-2.71309130e-12    2
 8.28515073e+04-3.29058903e+03-2.61093261e+02 3.59364993e+00-3.40538889e-03    3
 1.62077533e-06-3.02628703e-10 3.14263332e+05 1.20908943e+03                   4
BIN5BJ                                      G    300.00   3500.00 1390.00      1&
C 320.00 H 63.00 
 5.44961812e+02 5.40177677e-01-1.51289939e-04 1.27524221e-08 4.04609712e-13    2
-1.17297639e+05-2.91927429e+03-2.77265764e+02 2.90630020e+00-2.70465956e-03    3
 1.23739013e-06-2.19853971e-10 1.11281627e+05 1.31826109e+03                   4
BIN5CJ                                      G    300.00   3500.00 1370.00      1&
C 320.00 H 17.00 
 5.17964080e+02 4.57078766e-01-1.13727712e-04 4.66655739e-09 1.08851699e-12    2
-1.94746518e+05-2.88091788e+03-2.88688165e+02 2.81226780e+00-2.69240184e-03    3
 1.25949582e-06-2.27894924e-10 2.62761976e+04 1.26465571e+03                   4
BIN6AJ                                      G    300.00   3500.00 1290.00      1&
C 640.00 H 431.00 
 1.23762821e+03 1.77026241e+00-6.22545371e-04 9.54207658e-08-5.13173999e-12    2
 1.25536835e+05-6.67884001e+03-5.26755261e+02 7.24121890e+00-6.98412269e-03    3
 3.38305762e-06-6.42270665e-10 5.80747770e+05 2.28257683e+03                   4
BIN6BJ                                      G    300.00   3500.00 1390.00      1&
C 640.00 H 127.00 
 1.08992363e+03 1.08035536e+00-3.02579890e-04 2.55048499e-08 8.09218683e-13    2
-2.94595285e+05-5.83854863e+03-5.54531539e+02 5.81260044e+00-5.40931919e-03    3
 2.47478029e-06-4.39707947e-10 1.62563251e+05 2.63652221e+03                   4
BIN6CJ                                      G    300.00   3500.00 1370.00      1&
C 640.00 H 33.00 
 1.03577702e+03 9.08543668e-01-2.24434087e-04 8.57368301e-09 2.24989094e-12    2
-4.53333367e+05-5.76580457e+03-5.77679845e+02 5.61936664e+00-5.38226945e-03    3
 2.51846924e-06-4.55760247e-10-1.12461852e+04 2.52612570e+03                   4
BIN7AJ                                      G    300.00   3500.00 1260.00      1&
C 1250.00 H 812.00 
 2.35938249e+03 3.50442304e+00-1.25852280e-03 2.00397985e-07-1.15957197e-11    2
 2.45225502e+05-1.29759728e+04-1.05686227e+03 1.43496445e+01-1.41695007e-02    3
 7.03160324e-06-1.36699359e-09 1.10611918e+06 4.29496756e+03                   4
BIN7BJ                                      G    300.00   3500.00 1390.00      1&
C 1250.00 H 249.00 
 2.12942777e+03 2.10904362e+00-5.90181843e-04 4.95662128e-08 1.60771953e-12    2
-6.31142548e+05-1.14103717e+04-1.08227805e+03 1.13513625e+01-1.05639073e-02    3
 4.83312758e-06-8.58745044e-10 2.61711671e+05 5.14187909e+03                   4
BIN7CJ                                      G    300.00   3500.00 1370.00      1&
C 1250.00 H 64.00 
 2.02255555e+03 1.77107533e+00-4.36628637e-04 1.63379652e-08 4.43166058e-12    2
-9.45844123e+05-1.12606232e+04-1.12888932e+03 1.09723742e+01-1.05110435e-02    3
 4.91872961e-06-8.90165354e-10-8.23482304e+04 4.93538523e+03                   4
BIN8AJ                                      G    300.00   3500.00 1250.00      1&
C 2500.00 H 1562.00 
 4.78397135e+03 6.73406816e+00-2.34092722e-03 3.50725031e-07-1.79620968e-11    2
 4.78866181e+05-2.68188359e+04-2.11920594e+03 2.88242355e+01-2.88491280e-02    3
 1.44884321e-05-2.84550351e-09 2.20466050e+06 8.02540356e+03                   4
BIN8BJ                                      G    300.00   3500.00 1390.00      1&
C 2500.00 H 499.00 
 4.25751413e+03 4.22013813e+00-1.18195266e-03 9.96282958e-08 3.16101376e-12    2
-1.32524861e+06-2.28068302e+04-2.16613876e+03 2.27054702e+01-2.11301527e-02    3
 9.66711033e-06-1.71760914e-09 4.60526889e+05 1.02989147e+04                   4
BIN8CJ                                      G    300.00   3500.00 1370.00      1&
C 2500.00 H 125.00 
 4.04548911e+03 3.52987664e+00-8.66404388e-04 3.09041878e-08 9.03679946e-12    2
-1.95771333e+06-2.25361925e+04-2.25759576e+03 2.19330441e+01-2.10158578e-02    3
 9.83599103e-06-1.78021262e-09-2.30668072e+05 9.85682723e+03                   4
BIN9AJ                                      G    300.00   3500.00 1450.00      1&
C 5000.00 H 2999.00 
 9.86127424e+03 1.17426301e+01-3.79533336e-03 4.94630822e-07-1.77255210e-11    2
 5.82013094e+05-4.82475064e+04-3.84224391e+03 4.95454388e+01-4.29016872e-02    3
 1.84745636e-05-3.11771393e-09 4.55603336e+06 2.29557753e+04                   4
BIN9BJ                                      G    300.00   3500.00 1390.00      1&
C 5000.00 H 999.00 
 8.51502838e+03 8.44027594e+00-2.36390508e-03 1.99256525e-07 6.32203498e-12    2
-2.71049726e+06-4.56136613e+04-4.33227753e+03 4.54109404e+01-4.22603056e-02    3
 1.93342208e-05-3.43521830e-09 8.61053782e+05 2.05978292e+04                   4
BIN9CJ                                      G    300.00   3500.00 1370.00      1&
C 5000.00 H 250.00 
 8.09124297e+03 7.05642313e+00-1.73089314e-03 6.13022999e-08 1.81238981e-11    2
-3.97651917e+06-4.50778750e+04-4.51494854e+03 4.38628217e+01-4.20298697e-02    3
 1.96715099e-05-3.56038113e-09-5.22422694e+05 1.97082765e+04                   4
BIN10AJ                                     G    300.00   3500.00 1450.00      1&
C 10000.00 H 5749.00 
 1.97029151e+04 2.27863789e+01-7.21557544e-03 8.95246620e-07-2.64550359e-11    2
 6.35689932e+05-9.69907736e+04-7.72023177e+03 9.84364391e+01-8.54742584e-02    3
 3.68762503e-05-6.23007636e-09 8.58840251e+06 4.54994997e+04                   4
BIN10BJ                                     G    300.00   3500.00 1390.00      1&
C 10000.00 H 1999.00 
 1.70300565e+04 1.68805527e+01-4.72781083e-03 3.98513272e-07 1.26440433e-11    2
-5.48099451e+06-9.12273215e+04-8.66455517e+03 9.08218813e+01-8.45206115e-02    3
 3.86684417e-05-6.87043660e-09 1.66210755e+06 4.11956590e+04                   4
BIN10CJ                                     G    300.00   3500.00 1370.00      1&
C 10000.00 H 500.00 
 1.61813900e+04 1.41116083e+01-3.46149046e-03 1.22604030e-07 3.62425990e-11    2
-8.01708723e+06-9.01472220e+04-9.03123353e+03 8.77251076e+01-8.40602123e-02    3
 3.93433933e-05-7.12083573e-09-1.10882839e+06 3.94263168e+04                   4
BIN11AJ                                     G    300.00   3500.00 1440.00      1&
C 20000.00 H 10999.00 
 3.85320627e+04 4.57711908e+01-1.47699876e-02 1.91821759e-06-6.79480097e-11    2
 5.99191148e+05-1.90340584e+05-1.56381168e+04 1.96243912e+02-1.71512405e-01    3
 7.44841516e-05-1.26662004e-08 1.62002028e+07 9.07520012e+04                   4
BIN11BJ                                     G    300.00   3500.00 1390.00      1&
C 20000.00 H 3999.00 
 3.40601131e+04 3.37611051e+01-9.45562146e-03 7.97026463e-07 2.52880982e-11    2
-1.10219890e+07-1.82454643e+05-1.73291103e+04 1.81643762e+02-1.69041223e-01    3
 7.73368832e-05-1.37408732e-08 3.26421511e+06 8.23913177e+04                   4
BIN11CJ                                     G    300.00   3500.00 1370.00      1&
C 20000.00 H 1000.00 
 3.23630441e+04 2.82198873e+01-6.92106537e-03 2.44701921e-07 7.25355111e-11    2
-1.60952666e+07-1.80299930e+05-1.80622236e+04 1.75446946e+02-1.68118575e-01    3
 7.86863124e-05-1.42416270e-08-2.27874323e+06 7.88472539e+04                   4
BIN12AJ                                     G    300.00   3500.00 1430.00      1&
C 40000.00 H 20999.00 
 7.53518226e+04 9.18832287e+01-3.01846305e-02 4.08352367e-06-1.65200164e-10    2
-9.55187507e+04-3.73613199e+05-3.16727997e+04 3.91252802e+02-3.44208658e-01    3
 1.50481672e-04-2.57592820e-08 3.05135232e+07 1.80998711e+05                   4
BIN12BJ                                     G    300.00   3500.00 1390.00      1&
C 40000.00 H 7999.00 
 6.81202262e+04 6.75222092e+01-1.89112417e-02 1.59405249e-06 5.05762487e-11    2
-2.21039777e+07-3.64909286e+05-3.46582201e+04 3.63287522e+02-3.38082443e-01    3
 1.54673765e-04-2.74817462e-08 6.46843035e+06 1.64782634e+05                   4
BIN12CJ                                     G    300.00   3500.00 1370.00      1&
C 40000.00 H 2000.00 
 6.47263536e+04 5.64364445e+01-1.38402158e-02 4.88898133e-07 1.45121269e-10    2
-3.22516262e+07-3.60605353e+05-3.61242050e+04 3.50890630e+02-3.36235310e-01    3
 1.57372156e-04-2.84832104e-08-4.61857309e+06 1.57689135e+05                   4
BIN13AJ                                     G    300.00   3500.00 1430.00      1&
C 80000.00 H 39999.00 
 1.50544994e+05 1.78173818e+02-5.73666391e-02 7.41412093e-06-2.58322030e-10    2
-4.01088351e+06-7.51156625e+05-6.36406012e+04 7.77294363e+02-6.85814763e-01    3
 3.00396929e-04-5.14790927e-08 5.72461966e+07 3.58773772e+05                   4
BIN13BJ                                     G    300.00   3500.00 1390.00      1&
C 80000.00 H 15999.00 
 1.36240456e+05 1.35044414e+02-3.78224820e-02 3.18810499e-06 1.01152470e-10    2
-4.42679579e+07-7.29818595e+05-6.93164425e+04 7.26575057e+02-6.76164903e-01    3
 3.09347539e-04-5.49634940e-08 1.28768599e+07 3.29565274e+05                   4
BIN13CJ                                     G    300.00   3500.00 1370.00      1&
C 80000.00 H 4000.00 
 1.29452967e+05 1.12869565e+02-2.76785175e-02 9.77290080e-07 2.90292897e-10    2
-6.45643415e+07-7.21216164e+05-7.22481635e+04 7.01777975e+02-6.72468748e-01    3
 3.14743825e-04-5.69663741e-08-9.29823179e+06 3.15372879e+05                   4
BIN14AJ                                     G    300.00   3500.00 1420.00      1&
C 160000.00 H 75999.00 
 2.94370543e+05 3.57500522e+02-1.17188538e-01 1.57854625e-05-6.30992005e-10    2
-1.30784480e+07-1.47478168e+06-1.28888380e+05 1.54977918e+03-1.37663782e+00    3
 6.07076207e-04-1.04731475e-07 1.07127086e+08 7.15616609e+05                   4
BIN14BJ                                     G    300.00   3500.00 1390.00      1&
C 160000.00 H 31999.00 
 2.72480905e+05 2.70088841e+02-7.56449720e-02 6.37621196e-06 2.02304741e-10    2
-8.85959122e+07-1.45963715e+06-1.38632883e+05 1.45315010e+03-1.35232978e+00    3
 6.18695067e-04-1.09926986e-07 2.56937208e+07 6.59130542e+05                   4
BIN14CJ                                     G    300.00   3500.00 1370.00      1&
C 160000.00 H 8000.00 
 2.58906205e+05 2.25735790e+02-5.53551155e-02 1.95407343e-06 5.80636118e-10    2
-1.29189780e+08-1.44243786e+06-1.44496088e+05 1.40355270e+03-1.34493568e+00    3
 6.29487193e-04-1.13932707e-07-1.86575518e+07 6.30740392e+05                   4
BIN15AJ                                     G    300.00   3500.00 1420.00      1&
C 320000.00 H 143999.00 
 5.88112729e+05 6.92613672e+02-2.22352127e-01 2.85542667e-05-9.73083776e-10    2
-4.12583940e+07-2.96531673e+06-2.58962261e+05 3.07874040e+03-2.74290854e+00    3
 1.21191408e-03-2.09311080e-07 1.99310903e+08 1.41836311e+06                   4
BIN15BJ                                     G    300.00   3500.00 1390.00      1&
C 320000.00 H 63999.00 
 5.44961812e+05 5.40177677e+02-1.51289939e-01 1.27524221e-05 4.04609712e-10    2
-1.77251824e+08-2.91927429e+06-2.77265764e+05 2.90630020e+03-2.70465956e+00    3
 1.23739013e-03-2.19853971e-07 5.13274419e+07 1.31826109e+06                   4
BIN15CJ                                     G    300.00   3500.00 1370.00      1&
C 320000.00 H 16000.00 
 5.17812664e+05 4.51468257e+02-1.10708313e-01 3.90763869e-06 1.16132287e-09    2
-2.58440644e+08-2.88488114e+06-2.88991923e+05 2.80710209e+03-2.68986944e+00    3
 1.25897388e-03-2.27865364e-07-3.73761875e+07 1.26147536e+06                   4
BIN16AJ                                     G    300.00   3500.00 1410.00      1&
C 640000.00 H 271999.00 
 1.14984872e+06 1.38902743e+03-4.54050915e-01 6.08180693e-05-2.39260277e-09    2
-1.02799288e+08-5.82336592e+06-5.24438713e+05 6.13877902e+03-5.50697815e+00    3
 2.44990896e-03-4.25990278e-07 3.69349770e+08 2.82937106e+06                   4
BIN16BJ                                     G    300.00   3500.00 1390.00      1&
C 640000.00 H 127999.00 
 1.08992363e+06 1.08035536e+03-3.02579890e-01 2.55048499e-05 8.09218682e-10    2
-3.54563654e+08-5.83854863e+06-5.54531539e+05 5.81260044e+03-5.40931919e+00    3
 2.47478029e-03-4.39707947e-07 1.02594882e+08 2.63652221e+06                   4
BIN16CJ                                     G    300.00   3500.00 1370.00      1&
C 640000.00 H 32000.00 
 1.03562561e+06 9.02933158e+02-2.21414689e-01 7.81476413e-06 2.32269685e-09    2
-5.16942385e+08-5.76976784e+06-5.77983602e+05 5.61420092e+03-5.37973706e+00    3
 2.51794730e-03-4.55730686e-07-7.48134613e+07 2.52294535e+06                   4
BIN17AJ                                     G    300.00   3500.00 1410.00      1&
C 1250000.00 H 499999.00 
 2.24336632e+06 2.62543188e+03-8.39792285e-01 1.06983069e-04-3.54234720e-09    2
-2.59600475e+08-1.14354149e+07-1.02894704e+06 1.19085903e+04-1.07154928e+01    3
 4.77634500e-03-8.31443400e-07 6.63191892e+08 5.47593863e+06                   4
BIN17BJ                                     G    300.00   3500.00 1390.00      1&
C 1250000.00 H 249999.00 
 2.12875709e+06 2.11006902e+03-5.90976305e-01 4.98141439e-05 1.58050718e-09    2
-6.92564322e+08-1.14034153e+07-1.08306939e+06 1.13527352e+04-1.05650765e+01    3
 4.83355523e-03-8.58804580e-07 2.00323441e+08 5.14945736e+06                   4
BIN17CJ                                     G    300.00   3500.00 1370.00      1&
C 1250000.00 H 62500.00 
 2.02270654e+06 1.76353815e+03-4.32448787e-01 1.52627526e-05 4.53656195e-09    2
-1.00971136e+09-1.12690833e+07-1.12887404e+06 1.09652333e+04-1.05072975e+01    3
 4.91786552e-03-8.90098980e-07-1.46178276e+08 4.92762268e+06                   4
BIN18AJ                                     G    300.00   3500.00 1400.00      1&
C 2500000.00 H 937499.00 
 4.38558769e+06 5.26265421e+03-1.71431490e+00 2.28010293e-04-8.78779022e-09    2
-5.99143997e+08-2.24625968e+07-2.08368147e+06 2.37462804e+04-2.15182001e+01    3
 9.65843180e-03-1.69279163e-06 1.21225137e+09 1.09246167e+07                   4
BIN18BJ                                     G    300.00   3500.00 1390.00      1&
C 2500000.00 H 499999.00 
 4.25751413e+06 4.22013813e+03-1.18195266e+00 9.96282958e-05 3.16101376e-09    2
-1.38518861e+09-2.28068302e+07-2.16613876e+06 2.27054702e+04-2.11301527e+01    3
 9.66711033e-03-1.71760914e-06 4.00586889e+08 1.02989147e+07                   4
BIN18CJ                                     G    300.00   3500.00 1370.00      1&
C 2500000.00 H 125000.00 
 4.04541324e+06 3.52707308e+03-8.64895642e-01 3.05249772e-05 9.07317800e-09    2
-2.01948372e+09-2.25381712e+07-2.25774773e+06 2.19304628e+04-2.10145924e+01    3
 9.83573021e-03-1.78019785e-06-2.92417609e+08 9.85523968e+06                   4
BIN19AJ                                     G    300.00   3500.00 1400.00      1&
C 5000000.00 H 1749999.00 
 8.76152982e+06 1.01750298e+04-3.24032542e+00 4.08742172e-04-1.30444581e-08    2
-1.43342916e+09-4.51722315e+07-4.18606228e+06 4.71681501e+04-4.28758114e+01    3
 1.92827831e-02-3.38340892e-06 2.19189663e+09 2.16489213e+07                   4
BIN19BJ                                     G    300.00   3500.00 1390.00      1&
C 5000000.00 H 999999.00 
 8.51502838e+06 8.44027594e+03-2.36390508e+00 1.99256525e-04 6.32203499e-09    2
-2.77043726e+09-4.56136613e+07-4.33227753e+06 4.54109404e+04-4.22603056e+01    3
 1.93342208e-02-3.43521830e-06 8.01113782e+08 2.05978292e+07                   4
BIN19CJ                                     G    300.00   3500.00 1370.00      1&
C 5000000.00 H 250000.00 
 8.09082677e+06 7.05414290e+03-1.72978949e+00 6.10494994e-05 1.81463996e-08    2
-4.03902858e+09-4.50763483e+07-4.51549530e+06 4.38609227e+04-4.20291834e+01    3
 1.96714602e-02-3.56039569e-06-5.84896330e+08 1.97104742e+07                   4
BIN20AJ                                     G    300.00   3500.00 1400.00      1&
C 10000000.00 H 3249999.00 
 1.75037676e+07 1.96495036e+04-6.10404245e+00 7.22927555e-04-1.70266682e-08    2
-3.33708008e+09-9.08385330e+07-8.40952271e+06 9.36874759e+04-8.54304414e+01    3
 3.84974032e-02-6.76246876e-06 3.91864121e+09 4.28972163e+07                   4
BIN20BJ                                     G    300.00   3500.00 1390.00      1&
C 10000000.00 H 1999999.00 
 1.70300565e+07 1.68805527e+04-4.72781083e+00 3.98513272e-04 1.26440433e-08    2
-5.54093451e+09-9.12273215e+07-8.66455517e+06 9.08218813e+04-8.45206115e+01    3
 3.86684417e-02-6.87043660e-06 1.60216755e+09 4.11956590e+07                   4
BIN20CJ                                     G    300.00   3500.00 1370.00      1&
C 10000000.00 H 500000.00 
 1.61816539e+07 1.41082826e+04-3.45957729e+00 1.22098583e-04 3.62928372e-08    2
-8.07811834e+09-9.01527025e+07-9.03099053e+06 8.77218429e+04-8.40583660e+01    3
 3.93429203e-02-7.12079142e-06-1.16985377e+09 3.94209437e+07                   4
BIN21AJ                                     G    300.00   3500.00 1400.00      1&
C 20000000.00 H 5999999.00 
 3.49689534e+07 3.78978912e+04-1.14548658e+01 1.25674090e-03-1.59287835e-08    2
-7.61454482e+09-1.82665219e+08-1.68938425e+07 1.86077308e+05-1.70218527e+02    3
 7.68584842e-02-1.35162401e-05 6.90703802e+09 8.49931824e+07                   4
BIN21BJ                                     G    300.00   3500.00 1390.00      1&
C 20000000.00 H 3999999.00 
 3.40601131e+07 3.37611051e+04-9.45562146e+00 7.97026463e-04 2.52880982e-08    2
-1.10819290e+10-1.82454643e+08-1.73291103e+07 1.81643762e+05-1.69041223e+02    3
 7.73368832e-02-1.37408732e-05 3.20427511e+09 8.23913177e+07                   4
BIN21CJ                                     G    300.00   3500.00 1370.00      1&
C 20000000.00 H 1000000.00 
 3.23633082e+07 2.82165614e+04-6.91915227e+00 2.44196525e-04 7.25857410e-08    2
-1.61562978e+10-1.80305412e+08-1.80619808e+07 1.75443682e+05-1.68116730e+02    3
 7.86858401e-02-1.42415828e-05-2.33976861e+09 7.88418812e+07                   4
BIN22AJ                                     G    300.00   3500.00 1400.00      1&
C 40000000.00 H 11999999.00 
 6.99379048e+07 7.57957844e+04-2.29097321e+01 2.51348176e-03-3.18575436e-08    2
-1.52291484e+10-3.65330427e+08-3.37876835e+07 3.72154608e+05-3.40437043e+02    3
 1.53716963e-01-2.70324792e-05 1.38140163e+10 1.69986358e+08                   4
BIN22BJ                                     G    300.00   3500.00 1390.00      1&
C 40000000.00 H 7999999.00 
 6.81202262e+07 6.75222092e+04-1.89112417e+01 1.59405249e-03 5.05762487e-08    2
-2.21639177e+10-3.64909286e+08-3.46582201e+07 3.63287522e+05-3.38082443e+02    3
 1.54673765e-01-2.74817462e-05 6.40849035e+09 1.64782634e+08                   4
BIN22CJ                                     G    300.00   3500.00 1370.00      1&
C 40000000.00 H 2000000.00 
 6.47266172e+07 5.64331166e+04-1.38383016e+01 4.88392483e-04 1.45171524e-07    2
-3.23126582e+10-3.60610837e+08-3.61239618e+07 3.50887362e+05-3.36233460e+02    3
 1.57371681e-01-2.84831659e-05-4.67959957e+09 1.57683755e+08                   4
BIN23AJ                                     G    300.00   3500.00 1400.00      1&
C 80000000.00 H 23999999.00 
 1.39875812e+08 1.51591568e+05-4.58194656e+01 5.02696436e-03-6.37152148e-08    2
-3.04583586e+10-7.30660869e+08-6.75753698e+07 7.44309230e+05-6.80874104e+02    3
 3.07433935e-01-5.40649600e-05 2.76279723e+10 3.39972729e+08                   4
BIN23BJ                                     G    300.00   3500.00 1390.00      1&
C 80000000.00 H 15999999.00 
 1.36240456e+08 1.35044414e+05-3.78224820e+01 3.18810499e-03 1.01152470e-07    2
-4.43278979e+10-7.29818595e+08-6.93164425e+07 7.26575057e+05-6.76164903e+02    3
 3.09347539e-01-5.49634940e-05 1.28169199e+10 3.29565274e+08                   4
BIN23CJ                                     G    300.00   3500.00 1370.00      1&
C 80000000.00 H 4000000.00 
 1.29453233e+08 1.12866235e+05-2.76766023e+01 9.76784169e-04 2.90343180e-07    2
-6.46253736e+10-7.21221656e+08-7.22479214e+07 7.01774715e+05-6.72466909e+02    3
 3.14743357e-01-5.69663306e-05-9.35925732e+09 3.15367509e+08                   4
BIN24AJ                                     G    300.00   3500.00 1400.00      1&
C 160000000.00 H 47999999.00 
 2.79751621e+08 3.03183140e+05-9.16389324e+01 1.00539288e-02-1.27430401e-07    2
-6.09167755e+10-1.46132172e+09-1.35150738e+08 1.48861845e+06-1.36174819e+03    3
 6.14867863e-01-1.08129919e-04 5.52558850e+10 6.79945445e+08                   4
BIN24BJ                                     G    300.00   3500.00 1390.00      1&
C 160000000.00 H 31999999.00 
 2.72480905e+08 2.70088841e+05-7.56449720e+01 6.37621195e-03 2.02304742e-07    2
-8.86558522e+10-1.45963715e+09-1.38632883e+08 1.45315010e+06-1.35232978e+03    3
 6.18695067e-01-1.09926986e-04 2.56337808e+10 6.59130542e+08                   4
BIN24CJ                                     G    300.00   3500.00 1370.00      1&
C 160000000.00 H 8000000.00 
 2.58906469e+08 2.25732465e+05-5.53532045e+01 1.95356898e-03 5.80686219e-07    2
-1.29250811e+11-1.44244334e+09-1.44495846e+08 1.40354944e+06-1.34493384e+03    3
 6.29486724e-01-1.13932663e-04-1.87185769e+10 6.30735021e+08                   4
BIN25AJ                                     G    300.00   3500.00 1400.00      1&
C 320000000.00 H 95999999.00 
 5.59503241e+08 6.06366279e+05-1.83277863e+02 2.01078565e-02-2.54860672e-07    2
-1.21833610e+11-2.92264343e+09-2.70301474e+08 2.97723689e+06-2.72349638e+03    3
 1.22973572e+00-2.16259836e-04 1.10511711e+11 1.35989089e+09                   4
BIN25BJ                                     G    300.00   3500.00 1390.00      1&
C 320000000.00 H 63999999.00 
 5.44961812e+08 5.40177677e+05-1.51289939e+02 1.27524221e-02 4.04609712e-07    2
-1.77311764e+11-2.91927429e+09-2.77265764e+08 2.90630020e+06-2.70465956e+03    3
 1.23739013e+00-2.19853971e-04 5.12675019e+10 1.31826109e+09                   4
BIN25CJ                                     G    300.00   3500.00 1370.00      1&
C 320000000.00 H 16000000.00 
 5.17812933e+08 4.51464927e+05-1.10706401e+02 3.90713402e-03 1.16137298e-06    2
-2.58501678e+11-2.88488666e+09-2.88991684e+08 2.80709885e+06-2.68986762e+03    3
 1.25897342e+00-2.27865322e-04-3.74372131e+10 1.26147000e+09                   4
CSOLID                  C   1               G    300.00   3500.00 1500.00      1
 1.91389821e+00 8.92963112e-04-1.78036753e-07-1.58310714e-12 3.19362075e-15    2
-8.88852183e+02-1.10895704e+01-8.87506283e-01 8.36337508e-03-7.64844873e-06    3
 3.31859999e-09-5.50170229e-13-4.84308363e+01 3.56145864e+00                   4


! ---------------------------------------------------------------------------- !
! Thermodynamics from Lacroix et al. (2016)
! ---------------------------------------------------------------------------- !
C.(S)             J 3/67C   1H   0N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
H(S)              J 3/67C   0H   1N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
CH3(S)            J 3/67C   1H   3N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
C(B)              J 3/67C   1H   0N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
Ca(B)             J 3/67C   1H   0N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
CHCH.(S)          J 3/67C   2H   2N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
CH2CH2.(S)        J 3/67C   2H   4N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
CCH(S)            J 3/67C   2H   1N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
CH2CH2(S)         J 3/67C   2H   4N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
CH.CH2(S)         J 3/67C   2H   3N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
CHCH2(S)          J 3/67C   2H   3N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
C.CH2(S)          J 3/67C   2H   2N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
p1(S)             J 3/67C   3H   4N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
p2(S)             J 3/67C   3H   4N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
p3(S)             J 3/67C   3H   6N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
p3-2(S)           J 3/67C   3H   6N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
p4(S)             J 3/67C   3H   6N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
p5(S)             J 3/67C   3H   5N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
p6(S)             J 3/67C   3H   4N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
p6-2(S)           J 3/67C   3H   4N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
p7(S)             J 3/67C   3H   4N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
CH2CH3(S)         J 3/67C   2H   5N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
CH2.(S)           J 3/67C   1H   2N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
C6H6.(S)          J 3/67C   6H   6N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
C6H6(S)           J 3/67C   6H   6N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
C6H5.(S)          J 3/67C   6H   5N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
C6H5#(S)          J 3/67C   6H   5N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
c1(S)             J 3/67C   4H   8N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
c2(S)             J 3/67C   4H   8N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
c3(S)             J 3/67C   4H   8N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
c4(S)             J 3/67C   4H   7N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
c5(S)             J 3/67C   4H   6N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
c6(S)             J 3/67C   4H   6N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
c7(S)             J 3/67C   4H   6N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
c8(S)             J 3/67C   4H   5N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
c9(S)             J 3/67C   4H   4N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
c10(S)            J 3/67C   4H   4N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
c11(S)            J 3/67C   4H   4N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
c12(S)            J 3/67C   4H   3N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
c13(S)            J 3/67C   4H   4N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
c14(S)            J 3/67C   4H   4N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
C10H8.(1)(S)      J 3/67C  10H   8N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
C10H8(1)(S)       J 3/67C  10H   8N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
C10H7.(1)(S)      J 3/67C  10H   7N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
C10H8.(2)(S)      J 3/67C  10H   8N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
C10H8(2)(S)       J 3/67C  10H   8N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
C10H7.(2)(S)      J 3/67C  10H   7N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
CHC.(C6H5)(S)     J 3/67C   8H   6N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
C(C6H5)CH.(S)     J 3/67C   8H   6N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
CH.CH3(S)         J 3/67C   2H   4N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
CHCH2.(S)         J 3/67C   2H   3N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
C6H5C2H.1(S)      J 3/67C   8H   6N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
C6H5C2H.2(S)      J 3/67C   8H   6N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
C6H5C2H3.1(S)     J 3/67C   8H   8N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
C6H5C2H3.2(S)     J 3/67C   8H   8N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
C6H5C2H31(S)      J 3/67C   8H   8N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
C6H5C2H31-2.(S)   J 3/67C   8H   7N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
CH2CHCH.(S)       J 3/67C   3H   4N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
CH2CH2CH2.(S)     J 3/67C   3H   6N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
CHCH2cyc1(S)      J 3/67C   2H   3N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
CHCH.cyc1(S)      J 3/67C   2H   2N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
CHCH2cyc2(S)      J 3/67C   2H   3N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
CHCH.cyc2(S)      J 3/67C   2H   2N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
CH2CH2cyc1(S)     J 3/67C   2H   4N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
CH2CH.cyc1(S)     J 3/67C   2H   3N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
CH2c5(S)          J 3/67C   1H   2N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
CH.c5(S)          J 3/67C   1H   1N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
CHCH3c5(S)        J 3/67C   2H   4N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
C.CH3c5(S)        J 3/67C   2H   3N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
CH2CHCH.c5(S)     J 3/67C   3H   4N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
CHCH2CH2.Bz(S)    J 3/67C   3H   5N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
CHCH2CH2Bz(S)     J 3/67C   3H   5N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
Hz(S)             J 3/67C   0H   1N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
C.z(S)            J 3/67C   1H   0N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
CH3z(S)           J 3/67C   1H   3N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
CH2.z(S)          J 3/67C   1H   2N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
CH2CHCH.z(S)      J 3/67C   3H   4N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
CH2Bz(S)          J 3/67C   1H   2N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
CHCHz(S)          J 3/67C   2H   2N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
CHCHCH3z(S)       J 3/67C   3H   5N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
CHCHCH2.z(S)      J 3/67C   3H   4N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
CHCH.z(S)         J 3/67C   2H   2N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
CH.Bz(S)          J 3/67C   1H   1N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4 
CHCH3Bz(S)        J 3/67C   2H   4N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4 
CHCH2.Bz(S)       J 3/67C   2H   3N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4 
CH2CHz(S)         J 3/67C   2H   3N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4 
CH.CHz(S)         J 3/67C   2H   2N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4 
CH2CH2.z(S)       J 3/67C   2H   4N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4 
CH2CH2CH3z(S)     J 3/67C   3H   7N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4 
CH.CH2CH3z(S)     J 3/67C   3H   6N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4 
CH2CH2CH2.z(S)    J 3/67C   3H   6N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4 
CH2CH2z(S)        J 3/67C   2H   4N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4 
CH.CH2z(S)        J 3/67C   2H   3N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
CHC.z(S)          J 3/67C   2H   1N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4 
CHCCHCH.z(S)      J 3/67C   4H   3N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4 
CH2CH3z(S)        J 3/67C   2H   5N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4 
CH.CH3z(S)        J 3/67C   2H   4N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4 
CHCH2z(S)         J 3/67C   2H   3N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4 
CHCH2CH3Bz(S)     J 3/67C   3H   6N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4 
CHCH.CH3Bz(S)     J 3/67C   3H   5N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4 
CHCCH3Bz(S)       J 3/67C   3H   4N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4 
CHCCH2.Bz(S)      J 3/67C   3H   3N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4 
CHCHc5(S)         J 3/67C   2H   2N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4 
CHCc5(S)          J 3/67C   2H   1N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4 
CH2c5z(S)         J 3/67C   1H   2N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4 
CH.c5z(S)         J 3/67C   1H   1N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4 
CHCH3c5z(S)       J 3/67C   2H   4N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4 
C.CH3c5z(S)       J 3/67C   2H   3N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4 
CHCH2CH2c6z(S)    J 3/67C   3H   3N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4 
CHCH.CH2c6z(S)    J 3/67C   3H   3N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4 
CH2c5CHCH.z(S)    J 3/67C   3H   4N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
CH2c5z(S)         J 3/67C   1H   2N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
CHCHCHCH.z(S)     J 3/67C   4H   4N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
CH.CHCH2CHz(S)    J 3/67C   4H   5N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
CHCCHCHCHCH.z(S)  J 3/67C   6H   5N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
CH2CHCHCHCH.z(S)  J 3/67C   5H   6N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
C.CH3Bz(S)        J 3/67C   2H   3N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
CCH2Bz(S)         J 3/67C   2H   2N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
CCH.Bz(S)         J 3/67C   2H   1N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
CHC.CH3z(S)       J 3/67C   3H   4N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
CHC.z(S)          J 3/67C   2H   1N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
CHCCHCH.z(S)      J 3/67C   4H   3N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
CHCCH2CH2.z(S)    J 3/67C   4H   5N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
CCHCH3BZ(S)       J 3/67C   3H   4N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
CCHCH2.Bz(S)      J 3/67C   3H   3N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
CHC.z(S)          J 3/67C   3H   4N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
CHCCHCH.z(S)      J 3/67C   3H   4N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
CHCCH2CH2.z(S)    J 3/67C   3H   4N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
CHCCH3z(S)        J 3/67C   3H   4N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
CHCCH2.z(S)       J 3/67C   3H   3N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
CHCCH2c5z(S)      J 3/67C   3H   3N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
CHCCH2.z(S)       J 3/67C   3H   3N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
CHCCH.c5z(S)      J 3/67C   3H   2N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
CHCCHCH3c5z(S)    J 3/67C   4H   5N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
CHCC.CH3c5z(S)    J 3/67C   4H   4N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
CHCHCH.Bz(S)      J 3/67C   3H   3N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
CHCHCHBz(S)       J 3/67C   3H   3N   0     S   300.00   3000.00               1
 0.24753989E 01 0.88112187E-03-0.20939481E-06 0.42757187E-11 0.16006564E-13    2
-0.81255620E 03-0.12188747E 02 0.84197538E 00 0.83710416E-02-0.13077030E-04    3
 0.97593603E-08-0.27279380E-11-0.52486288E 03-0.45272678E 01                   4
styrene.1(S)            C   8H   8          G    300.00   4000.00 1000.00      1
 .157758892E+02 .965110900E-02-.942941600E-06-.546911100E-09 .102652200E-12    2
 .330269797E+05-.617628096E+02 .114355700E+00 .362732400E-01 .115828600E-05    3
-.219696400E-07 .846355600E-11 .383605400E+05 .238011700E+02                   4
styrene1(S)             C   8H   8          G    300.00   4000.00 1000.00      1
 .157758892E+02 .965110900E-02-.942941600E-06-.546911100E-09 .102652200E-12    2
 .330269797E+05-.617628096E+02 .114355700E+00 .362732400E-01 .115828600E-05    3
-.219696400E-07 .846355600E-11 .383605400E+05 .238011700E+02                   4
phenylac.1(S)           C   8H   6          G    300.00   4000.00 1000.00      1
 .157758892E+02 .965110900E-02-.942941600E-06-.546911100E-09 .102652200E-12    2
 .330269797E+05-.617628096E+02 .114355700E+00 .362732400E-01 .115828600E-05    3
-.219696400E-07 .846355600E-11 .383605400E+05 .238011700E+02                   4
C7H7(S)                 C   7H   7          S    200.00   3500.00 1600.00      1
 1.77148781e+01 1.72901839e-02-4.74309316e-06 3.88421745e-10 1.27959347e-14    2
 1.68881058e+04-7.24712964e+01-3.23806381e+00 6.96725387e-02-5.38515508e-05    3
 2.08502791e-08-3.18436927e-12 2.35930472e+04 3.84624951e+01                   4
C7H6.(S)                C   7H   6          G    300.00   3500.00 1290.00      1
 1.11282362e+01 2.73165807e-02-1.25329645e-05 2.76951413e-09-2.40721375e-13    2
 3.69620905e+04-3.50553513e+01-3.97785296e+00 7.41571673e-02-6.69987629e-05    3
 3.09172135e-08-5.69570188e-12 4.08594615e+04 4.16694449e+01                   4
 
END                                                       
