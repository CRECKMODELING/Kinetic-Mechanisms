! This thermodynamic database was obtained by fitting the thermodynamic properties
! extracted from the following file: thermo.CHEMKIN.CKT
! The thermodynamic properties are fitted in order to preserve not only the 
! continuity of each function at the intermediate temperature, but also the  continuity
! of the derivatives, from the 1st to the 3rd order
! The intermediate temperatures are chosen in order to minimize the fitting error.
! Last update: 11/20/2019

THERMO ALL
270.   1000.   3500.
!!!!!!!!!!!!!!!
!SOLID SPECIES!
!!!!!!!!!!!!!!!
CELL                    C   6H  10O   5     S 300.0    4000.0    1000.0        1
 2.92516210e+01 1.95010807e-02 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-1.25919988e+05 0.00000000e+00 2.92516210e+01 1.95010807e-02 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-1.25919988e+05 0.00000000e+00                   4
GMSW                    C   5H   8O   4     S 300.0    4000.0    1000.0        1
 2.38346742e+01 1.58897828e-02 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-1.03039895e+05 0.00000000e+00 2.38346742e+01 1.58897828e-02 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-1.03039895e+05 0.00000000e+00                   4
XYHW                    C   5H   8O   4     S 300.0    4000.0    1000.0        1
 2.38346742e+01 1.58897828e-02 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-1.07071125e+05 0.00000000e+00 2.38346742e+01 1.58897828e-02 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-1.07071125e+05 0.00000000e+00                   4
XYGR                    C   5H   8O   4     S 300.0    4000.0    1000.0        1
 2.38346742e+01 1.58897828e-02 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-1.09720219e+05 0.00000000e+00 2.38346742e+01 1.58897828e-02 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-1.09720219e+05 0.00000000e+00                   4
LIGC                    C  15H  14O   4     S 300.0    4000.0    1000.0        1
 4.65946547e+01 3.10631031e-02 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-1.03601488e+05 0.00000000e+00 4.65946547e+01 3.10631031e-02 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-1.03601488e+05 0.00000000e+00                   4
LIGH                    C  22H  28O   9     S 300.0    4000.0    1000.0        1
 7.87405700e+01 5.24937133e-02 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-2.24303494e+05 0.00000000e+00 7.87405700e+01 5.24937133e-02 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-2.24303494e+05 0.00000000e+00                   4
LIGO                    C  20H  22O  10     S 300.0    4000.0    1000.0        1
 7.62020414e+01 5.08013609e-02 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-2.51966073e+05 0.00000000e+00 7.62020414e+01 5.08013609e-02 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-2.51966073e+05 0.00000000e+00                   4
TGL                     C  57H 100O   7     S 300.0    4000.0    1000.0        1
 1.61902232e+02 1.07934821e-01 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-2.44625348e+05 0.00000000e+00 1.61902232e+02 1.07934821e-01 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-2.44625348e+05 0.00000000e+00                   4
TANN                    C  15H  12O   7     S 300.0    4000.0    1000.0        1
 5.48900197e+01 3.65933465e-02 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-1.59515809e+05 0.00000000e+00 5.48900197e+01 3.65933465e-02 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-1.59515809e+05 0.00000000e+00                   4
MOIST                   C   0H   2O   1     S 300.0    4000.0    1000.0        1   !From DH vaporization  engineering tool box
 9.04470000E+00 1.60000000E-03-6.00000000E-06 6.00000000E-09-2.00000000E-12    2
-3.70865499E+04-2.88280137E+02 9.04470000E+00 1.60000000E-03-6.00000000E-06    3
 6.00000000E-09-2.00000000E-12-3.70865499E+04-2.88280137E+02                   4
ASH                     C   0H   0K   1     S 300.0    4000.0    1000.0        1
 1.80625030E+01 1.20416687E-02 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
-1.55939610E+04 0.00000000E+00 1.80625030E+01 1.20416687E-02 0.00000000E+00    3
 0.00000000E+00	0.00000000E+00-1.55939610E+04 0.00000000E+00                   4
CELLA                   C   6H  10O   5     S 300.0    4000.0    1000.0        1
 2.92516210e+01 1.95010807e-02 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-1.25919988e+05 0.00000000e+00 2.92516210e+01 1.95010807e-02 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-1.25919988e+05 0.00000000e+00                   4
HCE1                    C   5H   8O   4     S 300.0    4000.0    1000.0        1
 2.38346742e+01 1.58897828e-02 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-9.92237373e+04 0.00000000e+00 2.38346742e+01 1.58897828e-02 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-9.92237373e+04 0.00000000e+00                   4
HCE2                    C   5H   8O   4     S 300.0    4000.0    1000.0        1
 2.38346742e+01 1.58897828e-02 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-1.10741538e+05 0.00000000e+00 2.38346742e+01 1.58897828e-02 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-1.10741538e+05 0.00000000e+00                   4
LIGCC                   C  15H  14O   4     S 300.0    4000.0    1000.0        1
 4.65946547e+01 3.10631031e-02 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-7.69910033e+04 0.00000000e+00 4.65946547e+01 3.10631031e-02 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-7.69910033e+04 0.00000000e+00                   4
LIGOH                   C  19H  22O   8     S 300.0    4000.0    1000.0        1
 6.82624420e+01 4.55082946e-02 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-1.86693370e+05 0.00000000e+00 6.82624420e+01 4.55082946e-02 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-1.86693370e+05 0.00000000e+00                   4
LIG                     C  11H  12O   4     S 300.0    4000.0    1000.0        1
 3.75634032e+01 2.50422688e-02 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-9.42255209e+04 0.00000000e+00 3.75634032e+01 2.50422688e-02 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-9.42255209e+04 0.00000000e+00                   4
ITANN                   C   8H   4O   4     S 300.0    4000.0    1000.0        1
 2.96079278e+01 1.97386186e-02 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-9.52526629e+04 0.00000000e+00 2.96079278e+01 1.97386186e-02 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-9.52526629e+04 0.00000000e+00                   4
CHAR                    C   1               S 300.0    4000.0    1000.0        1
-1.00796361E-01	4.99828606E-03 0.00000000E+00 0.00000000E+00 0.00000000E+00    2           
-1.94683964E+02 0.00000000E+00-1.00796361E-01 4.99828606E-03 0.00000000E+00    3
 0.00000000E+00	0.00000000E+00-1.94683964E+02 0.00000000E+00                   4 
CHARO                   C   1H   0O   1     S 300.0    4000.0    1000.0        1
-1.00796361E-01	4.99828606E-03 0.00000000E+00 0.00000000E+00 0.00000000E+00    2           
-1.94683964E+02 0.00000000E+00-1.00796361E-01 4.99828606E-03 0.00000000E+00    3
 0.00000000E+00	0.00000000E+00-1.94683964E+02 0.00000000E+00                   4 
COH2S                   C   1H   2O   1     S 300.0    4000.0    1000.0        1
 5.41694681e+00 3.61129787e-03 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-4.28130513e+04 0.00000000e+00 5.41694681e+00 3.61129787e-03 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-4.28130513e+04 0.00000000e+00                   4
CO2S                    C   1H   0O   2     S 300.0    4000.0    1000.0        1
 7.93959940e+00 5.29306627e-03 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-4.00155073e+04 0.00000000e+00 7.93959940e+00 5.29306627e-03 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-4.00155073e+04 0.00000000e+00                   4
COS                     C   1H   0O   1     S 300.0    4000.0    1000.0        1
 5.05324318e+00 3.36882879e-03 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-9.45019792e+03 0.00000000e+00 5.05324318e+00 3.36882879e-03 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-9.45019792e+03 0.00000000e+00                   4
COSTIFFS                C   1H   0O   1     S 300.0    4000.0    1000.0        1
 5.05324318e+00 3.36882879e-03 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-9.45019792e+03 0.00000000e+00 5.05324318e+00 3.36882879e-03 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-9.45019792e+03 0.00000000e+00                   4
CH3OHS                  C   1H   4O   1     S 300.0    4000.0    1000.0        1
 5.78065044e+00 3.85376696e-03 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-2.63330830e+04 0.00000000e+00 5.78065044e+00 3.85376696e-03 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-2.63330830e+04 0.00000000e+00                   4
CH4S                    C   1H   4O   0     S 300.0    4000.0    1000.0        1
 2.89429422e+00 1.92952948e-03 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-9.21591184e+03 0.00000000e+00 2.89429422e+00 1.92952948e-03 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-9.21591184e+03 0.00000000e+00                   4
C2H4S                   C   2H   4O   0     S 300.0    4000.0    1000.0        1
 5.06118118e+00 3.37412079e-03 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
 4.92120269e+03 0.00000000e+00 5.06118118e+00 3.37412079e-03 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00 4.92120269e+03 0.00000000e+00                   4
C6H5OHS                 C   6H   6O   1     S 300.0    4000.0    1000.0        1
 1.69787889e+01 1.13191926e-02 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-1.86144892e+04 0.00000000e+00 1.69787889e+01 1.13191926e-02 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-1.86144892e+04 0.00000000e+00                   4
CH2OS                   C   1H   2O   1     S 300.0    4000.0    1000.0        1
 5.41694681e+00 3.61129787e-03 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-2.45084187e+04 0.00000000e+00 5.41694681e+00 3.61129787e-03 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-2.45084187e+04 0.00000000e+00                   4
H2S                     C   0H   2O   0     S 300.0    4000.0    1000.0        1
 3.63703630e-01 2.42469087e-04 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
 1.09946128e+03 0.00000000e+00 3.63703630e-01 2.42469087e-04 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00 1.09946128e+03 0.00000000e+00                   4
C2H6S                   C   2H   6O   0     S 300.0    4000.0    1000.0        1
 5.42488481e+00 3.61658988e-03 0.00000000e+00 0.00000000e+00 0.00000000e+00    2
-1.10454007e+04 0.00000000e+00 5.42488481e+00 3.61658988e-03 0.00000000e+00    3
 0.00000000e+00 0.00000000e+00-1.10454007e+04 0.00000000e+00                   4

!!!!!!!!!!!!!
!GAS SPECIES!
!!!!!!!!!!!!! 

AR                      AR  1               G    200.00   3500.00  820.00      1
 2.50013930e+00-3.98275056e-07 3.45878291e-10-1.18292362e-13 1.38552083e-17    2
-7.45407890e+02 4.37897364e+00 2.49974490e+00 1.52564555e-06-3.17348868e-09    3
 2.74298160e-12-8.58484413e-16-7.45343208e+02 4.38079814e+00                   4
N2                      N   2               G    200.00   3500.00 1050.00      1
 2.81166076e+00 1.67067343e-03-6.79997337e-07 1.32881347e-10-1.02767403e-14    2
-8.69811587e+02 6.64838035e+00 3.73100682e+00-1.83159728e-03 4.32324654e-06    3
-3.04378144e-09 7.46071541e-13-1.06287426e+03 2.16821198e+00                   4
HE                      HE  1               G    200.00   3500.00  850.00      1
 2.50020615e+00-5.42574673e-07 4.63925536e-10-1.57302034e-13 1.82971341e-17    2
-7.45426807e+02 9.27648991e-01 2.49964853e+00 2.08151081e-06-4.16681355e-09    3
 3.47465019e-12-1.04992411e-15-7.45332012e+02 9.30248553e-01                   4
H2                      H   2               G    200.00   3500.00  700.00      1
 3.78199882e+00-1.01873257e-03 1.24226228e-06-4.19011878e-10 4.75543765e-14    2
-1.10283024e+03-5.60525913e+00 2.64204435e+00 5.49529297e-03-1.27163639e-05    3
 1.28749178e-08-4.70027765e-12-9.43236610e+02-5.12230966e-01                   4
H                       H   1               G    200.00   3500.00  860.00      1
 2.50031492e+00-7.73403020e-07 6.39349560e-10-2.12554687e-13 2.44483701e-17    2
 2.54736474e+04-4.48357210e-01 2.49950545e+00 2.99160564e-06-5.92752602e-09    3
 4.87804654e-12-1.45537757e-15 2.54737866e+04-4.44574039e-01                   4
O2                      O   2               G    200.00   3500.00  700.00      1
 2.82012407e+00 2.48211359e-03-1.51202095e-06 4.48556206e-10-4.87305673e-14    2
-9.31350151e+02 7.94914553e+00 3.74403921e+00-2.79740147e-03 9.80122559e-06    3
-1.03259643e-08 3.79931247e-12-1.06069827e+03 3.82132646e+00                   4
O                       O   1               G    200.00   3500.00  720.00      1
 2.62549144e+00-2.08959657e-04 1.33918551e-07-3.85875904e-11 4.38918689e-15    2
 2.92061519e+04 4.48358516e+00 3.14799200e+00-3.11174057e-03 6.18137878e-06    3
-5.63808780e-09 1.94866009e-12 2.91309118e+04 2.13446554e+00                   4
H2O                     H   2O   1          G    200.00   3500.00 1420.00      1
 2.66777069e+00 3.05768864e-03-9.00442530e-07 1.43361590e-10-1.00857860e-14    2
-2.98875645e+04 6.91191161e+00 4.06061172e+00-8.65807224e-04 3.24409535e-06    3
-1.80243084e-09 3.32483304e-13-3.02831314e+04-2.96150501e-01                   4
OH                      H   1O   1          G    200.00   3500.00 1700.00      1
 2.49867381e+00 1.66635254e-03-6.28251336e-07 1.28346754e-10-1.05735839e-14    2
 3.88110712e+03 7.78218797e+00 3.91354630e+00-1.66275921e-03 2.30920021e-06    3
-1.02359503e-09 1.58829619e-13 3.40005047e+03 2.05474752e-01                   4
H2O2                    H   2O   2          G    200.00   3500.00 1800.00      1
 4.76869611e+00 3.89237905e-03-1.21382388e-06 1.92615394e-10-1.22582099e-14    2
-1.80900219e+04-5.11810217e-01 3.34774226e+00 7.05005427e-03-3.84521989e-06    3
 1.16720651e-09-1.47618087e-13-1.75784785e+04 7.17868844e+00                   4
HO2                     H   1O   2          G    200.00   3500.00  700.00      1
 3.02391888e+00 4.46390908e-03-2.23146492e-06 6.12710797e-10-6.64266231e-14    2
 3.99341610e+02 9.10699976e+00 3.61994300e+00 1.05805693e-03 5.06678968e-06    3
-6.33800787e-09 2.41597290e-12 3.15898233e+02 6.44411476e+00                   4
CO                      C   1O   1          G    200.00   3500.00  960.00      1
 2.79255380e+00 1.87486885e-03-8.59711900e-07 1.91200058e-10-1.67855270e-14    2
-1.41723335e+04 7.41443564e+00 3.75723893e+00-2.14465251e-03 5.42079022e-06    3
-4.17025975e-09 1.11901130e-12-1.43575530e+04 2.79976793e+00                   4
CO2                     C   1O   2          G    200.00   3500.00 1450.00      1
 4.70876459e+00 2.62914723e-03-9.30606601e-07 1.43892961e-10-7.62581847e-15    2
-4.90562638e+04-2.34976404e+00 2.31684348e+00 9.22755029e-03-7.75654080e-06    3
 3.28225351e-09-5.48722465e-13-4.83626067e+04 1.00786234e+01                   4
HOCO                    H   1C   1O   2     G    200.00   3500.00 1570.00      1
 5.88810551e+00 3.28985483e-03-9.88703679e-07 1.12295220e-10-2.32818091e-15    2
-2.40914384e+04-5.05613781e+00 2.36661498e+00 1.22618052e-02-9.56063081e-06    3
 3.75217935e-09-5.81927565e-13-2.29856904e+04 1.35214769e+01                   4
CH4                     C   1H   4          G    300.00   3500.00  700.00      1
 5.05346544e-01 1.23697842e-02-4.99807893e-06 1.04392755e-09-8.62897300e-14    2
-9.58982509e+03 1.61752768e+01 5.23967275e+00-1.46835084e-02 5.29732624e-05    3
-5.41668737e-08 1.96318536e-11-1.02526308e+04-4.97649490e+00                   4
CH3                     C   1H   3          G    300.00   3500.00 1060.00      1
 2.78805103e+00 6.15233479e-03-2.21179351e-06 3.74402654e-10-2.48151355e-14    2
 1.65862829e+04 5.77899820e+00 3.47829310e+00 3.54764774e-03 1.47408440e-06    3
-1.94375955e-09 5.21921234e-13 1.64399516e+04 2.40875956e+00                   4
CH2                     C   1H   2          G    300.00   3500.00 1800.00      1
 2.81272979e+00 3.55431373e-03-1.28768512e-06 2.21273711e-10-1.48738112e-14    2
 4.62073492e+04 6.64284613e+00 3.76489460e+00 1.43839193e-03 4.75583051e-07    3
-4.31788574e-10 7.58292840e-14 4.58645699e+04 1.48953154e+00                   4
CH2(S)                  C   1H   2          G    300.00   3500.00  970.00      1
 2.75934299e+00 3.65468308e-03-1.35589915e-06 2.74980416e-10-2.36795479e-14    2
 5.06429079e+04 6.11646385e+00 4.18185434e+00-2.21134310e-03 7.71527536e-06    3
-5.95950379e-09 1.58314628e-12 5.03669407e+04-7.03002562e-01                   4
C                       C   1               G    200.00   3500.00  700.00      1
 2.49472530e+00 3.92839623e-05-6.70015037e-08 3.71818699e-11-5.07306880e-15    2
 8.54504422e+04 4.79314257e+00 2.54495193e+00-2.47725357e-04 5.48018467e-07    3
-5.48551435e-10 2.04117397e-13 8.54434105e+04 4.56874269e+00                   4
CH                      C   1H   1          G    300.00   3500.00 1590.00      1
 2.27990133e+00 2.16985229e-03-7.07637823e-07 1.23973477e-10-9.56348334e-15    2
 7.11059412e+04 8.77326037e+00 3.77264331e+00-1.58547346e-03 2.83512232e-06    3
-1.36146054e-09 2.23995325e-13 7.06312492e+04 8.79407939e-01                   4
CH3O2H                  C   1H   4O   2     G    300.00   3500.00 1090.00      1
 7.33435504e+00 9.33238581e-03-3.40995754e-06 5.79327833e-10-3.79241273e-14    2
-1.81046373e+04-1.19553967e+01 7.70006816e-01 3.34217371e-02-3.65604409e-05    3
 2.08548529e-08-4.68827390e-12-1.66736094e+04 2.02794894e+01                   4
CH3O2                   C   1H   3O   2     G    300.00   3500.00 1800.00      1
 5.64141552e+00 8.74328811e-03-3.21961767e-06 5.43696238e-10-3.45016043e-14    2
-1.19010046e+03-3.41913229e+00 1.44289655e+00 1.80733303e-02-1.09946528e-05    3
 3.42333889e-09-4.34451972e-13 3.21366368e+02 1.93041283e+01                   4
CH3OH                   C   1H   4O   1     G    300.00   3500.00 1800.00      1
 2.71701641e+00 1.21538330e-02-5.02106867e-06 1.01068022e-09-8.18460330e-14    2
-2.57693414e+04 9.47419935e+00 8.47330413e-01 1.63086907e-02-8.48345015e-06    3
 2.29304373e-09-2.59952076e-13-2.50962544e+04 1.95933300e+01                   4
CH3O                    C   1H   3O   1     G    300.00   3500.00 1740.00      1
 5.72237859e+00 5.90228063e-03-1.80341022e-06 2.13335899e-10-5.61825765e-15    2
-7.86244706e+01-7.49172569e+00 8.89661124e-01 1.70119760e-02-1.13807338e-05    3
 3.88280853e-09-5.32841337e-13 1.60316121e+03 1.85001128e+01                   4
CH2OH                   C   1H   3O   1     G    300.00   3500.00 1360.00      1
 5.04534911e+00 6.02727160e-03-2.11386901e-06 3.36086164e-10-2.00987773e-14    2
-4.03584131e+03-1.57523866e+00 2.34821584e+00 1.39600165e-02-1.08632200e-05    3
 4.62498372e-09-8.08499063e-13-3.30222106e+03 1.22661975e+01                   4
CH2O                    C   1H   2O   1     G    300.00   3500.00  700.00      1
 1.33335656e+00 1.00905181e-02-5.12952546e-06 1.25425201e-09-1.19639101e-13    2
-1.39080170e+04 1.59916142e+01 4.32621275e+00-7.01151723e-03 3.15176932e-05    3
-3.36478610e-08 1.23454012e-11-1.43270169e+04 2.62028992e+00                   4
HCO                     C   1H   1O   1     G    200.00   3500.00  770.00      1
 2.60049318e+00 5.29278252e-03-2.69184204e-06 7.21357770e-10-7.43521372e-14    2
 4.05725330e+03 1.07450933e+01 4.03483982e+00-2.15836886e-03 1.18233879e-05    3
-1.18459409e-08 4.00593964e-12 3.83636392e+03 4.20008756e+00                   4
HO2CHO                  C   1H   2O   3     G    300.00   3500.00 1750.00      1
 1.00230822e+01 4.43559546e-03-1.56185376e-06 2.43414079e-10-1.38379679e-14    2
-3.81313379e+04-2.33591538e+01 2.47434347e+00 2.16898554e-02-1.63512194e-05    3
 5.87745813e-09-8.18701404e-13-3.54892793e+04 1.72835403e+01                   4
HOCHO                   H   2C   1O   2     G    200.00   3500.00 1800.00      1
 3.79473623e+00 8.42765802e-03-3.84722303e-06 8.63389995e-10-7.73674578e-14    2
-4.73118220e+04 5.12934093e+00 1.85206267e+00 1.27447104e-02-7.44476667e-06    3
 2.19581357e-09-2.62426287e-13-4.66124595e+04 1.56434955e+01                   4
OCHO                    C   1O   2H   1     G    200.00   3500.00  700.00      1
 2.58373953e+00 8.99565936e-03-4.55939784e-06 1.11902582e-09-1.07899897e-13    2
-1.67164582e+04 1.34890938e+01 4.25809176e+00-5.72067675e-04 1.59428744e-05    3
-1.84069477e-08 6.86566208e-12-1.69508675e+04 6.00851165e+00                   4
C2H6                    C   2H   6          G    300.00   3500.00 1800.00      1
 4.07959174e+00 1.57445255e-02-5.96197340e-06 1.06867166e-09-7.61012177e-14    2
-1.25948055e+04-1.43089592e+00-2.41778736e-01 2.53475710e-02-1.39645113e-05    3
 4.03257459e-09-4.87754402e-13-1.10391121e+04 2.19572626e+01                   4
C2H5                    C   2H   5          G    300.00   3500.00 1800.00      1
 5.19791696e+00 1.11042732e-02-3.71281218e-06 5.47664237e-10-2.89411242e-14    2
 1.17176203e+04-4.91384359e+00 6.75421537e-01 2.11542630e-02-1.20878037e-05    3
 3.64951295e-09-4.59753446e-13 1.33457186e+04 1.95628451e+01                   4
C2H5O2H                 C   2H   6O   2     G    300.00   3500.00 1450.00      1
 1.00876754e+01 1.40221795e-02-4.79127924e-06 7.15473842e-10-3.78163306e-14    2
-2.40669300e+04-2.56733607e+01-5.77204966e-01 4.34425392e-02-3.52261341e-05    3
 1.47085106e-08-2.45040887e-12-2.09741147e+04 2.97412033e+01                   4
C2H5O2                  C   2H   5O   2     G    300.00   3500.00 1480.00      1
 9.29919856e+00 1.29334585e-02-4.54028293e-06 7.01326950e-10-3.92077242e-14    2
-7.64002502e+03-2.14311828e+01 2.00183001e-01 3.75253925e-02-2.94645403e-05    3
 1.19284699e-08-1.93568458e-12-4.94671641e+03 2.60335046e+01                   4
C2H4                    C   2H   4          G    300.00   3500.00 1650.00      1
 4.60402750e+00 9.50595291e-03-3.15129224e-06 4.53051970e-10-2.23949056e-14    2
 3.97229090e+03-3.77421075e+00-6.02932966e-02 2.08133973e-02-1.34307871e-05    3
 4.60638323e-09-6.51687520e-13 5.51151677e+03 2.10642174e+01                   4
C2H3                    C   2H   3          G    300.00   3500.00 1450.00      1
 4.18728262e+00 7.47581866e-03-2.58984442e-06 4.05266469e-10-2.35023462e-14    2
 3.38403788e+04 1.51959352e+00 1.23421228e+00 1.56222196e-02-1.10171557e-05    3
 4.27989236e-09-6.91541292e-13 3.46967692e+04 1.68637042e+01                   4
C2H2                    C   2H   2          G    300.00   3500.00  790.00      1
 4.37267451e+00 5.47212841e-03-2.03181554e-06 3.75019163e-10-2.77049120e-14    2
 2.58626598e+04-2.43835909e+00 7.70536924e-01 2.37107997e-02-3.66622041e-05    3
 2.95989758e-08-9.27579245e-12 2.64317975e+04 1.40907683e+01                   4
C2H                     C   2H   1          G    300.00   3500.00 1710.00      1
 3.41788259e+00 4.21328984e-03-1.58936942e-06 2.68739179e-10-1.73346344e-14    2
 6.72874491e+04 5.32512356e+00 4.60873599e+00 1.42766785e-03 8.54158644e-07    3
-6.83903342e-10 1.21940588e-13 6.68801772e+04-1.05894068e+00                   4
C2H5OH                  C   2H   6O   1     G    300.00   3500.00 1580.00      1
 7.32490792e+00 1.39762984e-02-4.67366801e-06 6.82063840e-10-3.47025203e-14    2
-3.18909573e+04-1.38313053e+01-4.22291371e-01 3.35894612e-02-2.32937592e-05    3
 8.53864242e-09-1.27783204e-12-2.94428423e+04 2.70882144e+01                   4
C2H5O                   C   2H   5O   1     G    300.00   3500.00  700.00      1
 1.68957251e+00 2.35453826e-02-1.23415273e-05 3.08911892e-09-2.98016647e-13    2
-3.10347953e+03 1.69410915e+01 3.27852963e+00 1.44656276e-02 7.11509041e-06    3
-1.54409932e-08 6.31988055e-12-3.32593352e+03 9.84203310e+00                   4
PC2H4OH                 C   2H   5O   1     G    300.00   3500.00 1470.00      1
 7.18479728e+00 1.17471688e-02-4.06239662e-06 6.31554442e-10-3.61644761e-14    2
-6.24418465e+03-9.60110342e+00 1.82077783e+00 2.63431401e-02-1.89562449e-05    3
 7.38613415e-09-1.18490252e-12-4.66716293e+03 1.83437447e+01                   4
SC2H4OH                 C   2H   5O   1     G    300.00   3500.00 1500.00      1
 6.63757447e+00 1.19924580e-02-4.07718691e-06 6.22004854e-10-3.47507928e-14    2
-9.66525362e+03-7.65007915e+00 1.23305390e+00 2.64045128e-02-1.84892418e-05    3
 7.02736257e-09-1.10231041e-12-8.04389745e+03 2.06149530e+01                   4
C2H4O2H                 C   2H   5O   2     G    300.00   3500.00 1440.00      1
 9.66417590e+00 1.29483241e-02-4.44318413e-06 6.83406719e-10-3.84804652e-14    2
 1.86599146e+03-2.38806219e+01 2.23212425e+00 3.35929120e-02-2.59479632e-05    3
 1.06393230e-08-1.76693815e-12 4.00642233e+03 1.46847777e+01                   4
C2H4O1-2                C   2H   4O   1     G    300.00   3500.00 1520.00      1
 6.04215722e+00 1.11433665e-02-3.80167598e-06 5.65227352e-10-2.94248630e-14    2
-9.44151496e+03-1.02352874e+01-2.19672845e+00 3.28246446e-02-2.51976741e-05    3
 9.94943705e-09-1.57288040e-12-6.93689372e+03 3.29622800e+01                   4
C2H3O1-2                C   2H   3O   1     G    200.00   3500.00 1800.00      1
 7.60993641e+00 6.11300571e-03-1.59366922e-06 1.28294122e-10 2.98968411e-15    2
 1.61313301e+04-1.70584536e+01 7.34197611e-02 2.28608205e-02-1.55501815e-05    3
 5.29737275e-09-7.14937904e-13 1.88444761e+04 2.37307467e+01                   4
CH3CHO                  C   2H   4O   1     G    300.00   3500.00 1800.00      1
 6.22195717e+00 1.06589200e-02-3.75189849e-06 6.00730261e-10-3.66602428e-14    2
-2.30621368e+04-8.31410467e+00 9.75916365e-01 2.23167884e-02-1.34667889e-05    3
 4.19883781e-09-5.36397402e-13-2.11735621e+04 2.00785625e+01                   4
CH3CO                   C   2H   3O   1     G    300.00   3500.00 1800.00      1
 6.07689133e+00 8.12979100e-03-2.81854834e-06 4.38697836e-10-2.55171354e-14    2
-4.06801092e+03-6.15493095e+00 1.47388055e+00 1.83587038e-02-1.13426424e-05    3
 3.59576970e-09-4.63999338e-13-2.41092704e+03 1.87575236e+01                   4
CH2CHO                  C   2H   3O   1     G    300.00   3500.00 1340.00      1
 6.47703838e+00 7.91358487e-03-2.83605797e-06 4.62112353e-10-2.83230958e-14    2
-1.16170826e+03-8.37157531e+00 7.37868219e-01 2.50454361e-02-2.20135034e-05    3
 1.00031300e-08-1.80836370e-12 3.76389344e+02 2.09962839e+01                   4
CH2CO                   C   2H   2O   1     G    300.00   3500.00 1360.00      1
 5.69523630e+00 6.46841649e-03-2.33588407e-06 3.83408083e-10-2.36897816e-14    2
-8.05944305e+03-4.61154409e+00 2.49503978e+00 1.58807592e-02-1.27171444e-05    3
 5.47226118e-09-9.59140719e-13-7.18898960e+03 1.18115657e+01                   4
HCCO                    C   2H   1O   1     G    300.00   3500.00 1220.00      1
 5.81420551e+00 3.89116666e-03-1.41168512e-06 2.35668209e-10-1.49424599e-14    2
 1.94026781e+04-4.94089845e+00 3.33028657e+00 1.20351632e-02-1.14247956e-05    3
 5.70731328e-09-1.13618120e-12 2.00087543e+04 7.53650401e+00                   4
CH3CO3                  C   2H   3O   3     G    300.00   3500.00 1760.00      1
 1.40469371e+01 2.48483616e-03 1.65900305e-06-8.55133607e-10 9.82286856e-14    2
-2.73756812e+04-4.36816920e+01 2.64892556e+00 2.83894079e-02-2.04187569e-05    3
 7.50765427e-09-1.08966732e-12-2.33635811e+04 1.77505784e+01                   4
CH3CO3H                 C   2H   4O   3     G    300.00   3500.00 1240.00      1
 1.23807020e+01 1.08772141e-02-4.04888352e-06 6.94756538e-10-4.56573485e-14    2
-7.51809422e+04-3.74730284e+01-2.33886891e+00 5.83597007e-02-6.14873754e-05    3
 3.15756662e-08-6.27164719e-12-7.15304886e+04 3.67067395e+01                   4
CH2OHCHO                C   2H   4O   2     G    300.00   3500.00 1800.00      1
 8.91045191e+00 9.14305835e-03-2.53718679e-06 2.39203927e-10 8.50817753e-16    2
-4.09945451e+04-1.84179625e+01 1.56305394e+00 2.54706094e-02-1.61434793e-05    3
 5.27857153e-09-6.99061350e-13-3.83494818e+04 2.13476881e+01                   4
CHOCHO                  C   2H   2O   2     G    300.00   3500.00 1570.00      1
 9.97760190e+00 4.26981387e-03-1.12729558e-06 7.37812974e-11 5.98356282e-15    2
-2.96900175e+04-2.75230936e+01 7.08345804e-01 2.78857530e-02-2.36902947e-05    3
 9.65467265e-09-1.51963608e-12-2.67794711e+04 2.13768443e+01                   4
O2C2H4O2H               C   2H   5O   4     G    300.00   3500.00 1800.00      1
 1.24323233e+01 1.62358946e-02-6.84260441e-06 1.39267464e-09-1.12911160e-13    2
-1.87641101e+04-2.90906711e+01 5.81911533e+00 3.09319123e-02-1.90892858e-05    3
 5.92848256e-09-7.42884481e-13-1.63833552e+04 6.70138985e+00                   4
HO2CH2CHO               C   2H   4O   3     G    300.00   3500.00 1240.00      1
 1.23807020e+01 1.08772141e-02-4.04888352e-06 6.94756538e-10-4.56573485e-14    2
-7.51809422e+04-3.74730284e+01-2.33886891e+00 5.83597007e-02-6.14873754e-05    3
 3.15756662e-08-6.27164719e-12-7.15304886e+04 3.67067395e+01                   4
CH3OCHO                 C   2H   4O   2     G    300.00   3500.00  700.00      1
 5.02910653e+00-2.87377518e-02 6.15808969e-05-2.98073517e-08 4.29774801e-12    2
-4.07046731e+04 1.82412183e+01 3.04007016e-07-1.95406361e-09 4.40443198e-12    3
 2.88411173e-08-1.66481338e-11-4.00005982e+04 4.07099926e+01                   4
CH3OCO                  C   2H   3O   2     G    300.00   3500.00  730.00      1
 2.57527322e+00 2.11166692e-02-1.20149822e-05 3.14849391e-09-3.11411023e-13    2
-2.07588781e+04 1.60124233e+01 4.66126873e+00 9.68655681e-03 1.14715501e-05    3
-1.83003940e-08 7.03409854e-12-2.10634335e+04 6.60518603e+00                   4
C3H8                    C   3H   8          G    300.00   3500.00 1690.00      1
 8.33847138e+00 1.79340895e-02-5.80534794e-06 7.91037165e-10-3.43400666e-14    2
-1.70816238e+04-2.27461869e+01-1.38651279e+00 4.09518035e-02-2.62352716e-05    3
 8.85017865e-09-1.22652076e-12-1.37945792e+04 2.92742167e+01                   4
IC3H7                   C   3H   7          G    300.00   3500.00 1800.00      1
 6.05951179e+00 1.82035635e-02-6.54041412e-06 1.09272169e-09-7.13189609e-14    2
 7.29671845e+03-6.80792692e+00-6.08211152e-01 3.30207256e-02-1.88880492e-05    3
 5.66591987e-09-7.06485374e-13 9.69709871e+03 2.92791806e+01                   4
NC3H7                   C   3H   7          G    300.00   3500.00 1590.00      1
 7.21724942e+00 1.65877274e-02-5.58902508e-06 8.31338728e-10-4.40999556e-14    2
 8.50975649e+03-1.26938745e+01-1.37086151e-01 3.50892006e-02-2.30432450e-05    3
 8.14966994e-09-1.19478096e-12 1.08484352e+04 2.61969990e+01                   4
C3H6                    C   3H   6          G    298.00   3500.00 1800.00      1
 6.31755560e+00 1.65819945e-02-6.59971811e-06 1.29512777e-09-1.03784233e-13    2
-3.79457444e+02-1.05616384e+01-8.55990160e-02 3.08112270e-02-1.84574118e-05    3
 5.68686619e-09-7.13747903e-13 1.92567822e+03 2.40935701e+01                   4
C3H5-A                  C   3H   5          G    298.00   3500.00 1600.00      1
 8.53877816e+00 1.04611881e-02-3.15379681e-06 3.85306812e-10-1.26413619e-14    2
 1.71766363e+04-2.28181771e+01-3.57888141e-01 3.27028538e-02-2.40053585e-05    3
 9.07345750e-09-1.37016491e-12 2.00235695e+04 2.42845605e+01                   4
C3H5-S                  C   3H   5          G    300.00   3500.00 1800.00      1
 6.52599586e+00 1.37686641e-02-5.50691249e-06 1.07278340e-09-8.39559751e-14    2
 2.86430047e+04-9.99636084e+00 1.54227615e+00 2.48435968e-02-1.47360231e-05    3
 4.49097250e-09-5.58704461e-13 3.04371438e+04 1.69765699e+01                   4
C3H5-T                  C   3H   5          G    300.00   3500.00  770.00      1
 1.49331934e+00 2.33788729e-02-1.18550710e-05 2.86552468e-09-2.68203788e-13    2
 2.87117776e+04 1.76892214e+01 2.52238876e+00 1.80330577e-02-1.44114539e-06    3
-6.15086111e-09 2.65919419e-12 2.85533009e+04 1.29935189e+01                   4
C3H5O                   C   3H   5O   1     G    300.00   3500.00 1610.00      1
 9.11079932e+00 1.37589671e-02-5.15319282e-06 9.32422242e-10-6.74696193e-14    2
 7.77376182e+03-2.10036633e+01 9.27196877e-01 3.40908986e-02-2.40959862e-05    3
 8.77622901e-09-1.28545204e-12 1.04088818e+04 2.23747991e+01                   4
C3H6O                   C   3H   6O   1     G    300.00   3500.00 1550.00      1
 9.00938188e+00 1.57632599e-02-5.29374429e-06 7.64253653e-10-3.74126701e-14    2
-1.56669514e+04-2.44960160e+01-1.88321637e+00 4.38731909e-02-3.24969033e-05    3
 1.24645371e-08-1.92455516e-12-1.22902459e+04 3.28282089e+01                   4
CH3CHCHO                C   3H   5O   1     G    300.00   3500.00 1800.00      1
 6.70347438e+00 1.89922304e-02-9.18109881e-06 2.14445631e-09-1.96154611e-13    2
-6.21094393e+03-1.05801373e+01 2.92067419e-01 3.32398014e-02-2.10540747e-05    3
 6.54185478e-09-8.06904398e-13-3.90283742e+03 2.41197347e+01                   4
AC4H7OOH                C   4H   8O   2     G    300.00   3500.00 1660.00      1
 1.22738315e+01 2.55483291e-02-9.81264424e-06 1.82078478e-09-1.35039680e-13    2
-1.24525975e+04-3.36837710e+01 1.60151398e+00 5.12647569e-02-3.30503802e-05    3
 1.11532089e-08-1.54052523e-12-8.90938812e+03 2.32129103e+01                   4
CH3CHCO                 C   3H   4O   1     G    300.00   3500.00 1280.00      1
 6.99681438e+00 1.49445090e-02-6.71568613e-06 1.45955089e-09-1.25293211e-13    2
-1.29366479e+04-1.07908045e+01 1.50068785e+00 3.21199044e-02-2.68431026e-05    3
 1.19425803e-08-2.17275989e-12-1.15296395e+04 1.70816031e+01                   4
AC3H5OOH                C   3H   6O   2     G    298.00   3500.00 1800.00      1
 1.36957660e+01 1.27112955e-02-4.21186204e-06 6.49029927e-10-3.94931006e-14    2
-1.11479409e+04-4.31791036e+01 4.22354617e+00 3.37606729e-02-2.17530099e-05    3
 7.14575135e-09-9.41815521e-13-7.73794171e+03 8.08652620e+00                   4
C3H6OH1-2               C   3H   7O   1     G    300.00   3500.00 1800.00      1
 8.46016309e+00 1.89669011e-02-7.38013611e-06 1.39189593e-09-1.05413410e-13    2
-1.21581705e+04-1.51603301e+01 4.08605516e-01 3.68592513e-02-2.22904279e-05    3
 6.91422623e-09-8.72403729e-13-9.25960980e+03 2.84163791e+01                   4
C3H6OH2-1               C   3H   7O   1     G    300.00   3500.00 1590.00      1
 8.99548175e+00 1.75103805e-02-6.94615452e-06 1.37004351e-09-1.07539367e-13    2
-1.65436317e+04-1.93287204e+01 1.31207700e+00 3.68397006e-02-2.51813622e-05    3
 9.01583289e-09-1.30970751e-12-1.41003090e+04 2.13023222e+01                   4
HOC3H6O2                C   3H   7O   3     G    300.00   3500.00 1480.00      1
 1.24409054e+01 2.15172911e-02-8.97737608e-06 1.82414695e-09-1.48047126e-13    2
-3.10315628e+04-3.23089021e+01 2.93449050e+00 4.72103043e-02-3.50175922e-05    3
 1.35539740e-08-2.12943683e-12-2.82176640e+04 1.72809692e+01                   4
SC3H5OH                 C   3H   6O   1     G    300.00   3500.00 1260.00      1
 7.83167551e+00 1.85990423e-02-7.98421803e-06 1.67672179e-09-1.40411927e-13    2
-2.22362405e+04-1.56369779e+01-5.71229119e-02 4.36428468e-02-3.77982710e-05    3
 1.74513530e-08-3.27029907e-12-2.02482633e+04 2.42451081e+01                   4
C3H5OH                  C   3H   6O   1     G    300.00   3500.00 1630.00      1
 9.39463141e+00 1.51343100e-02-4.86246233e-06 6.64177119e-10-2.94552392e-14    2
-2.20582200e+04-2.45922041e+01 4.73537639e-01 3.70265647e-02-2.50087089e-05    3
 8.90395079e-09-1.29322421e-12-1.91499434e+04 2.28055846e+01                   4
CH2CCH2OH               C   3H   5O   1     G    300.00   3500.00 1800.00      1
 7.15397445e+00 1.62590917e-02-7.06959863e-06 1.52062077e-09-1.30983718e-13    2
 1.01359979e+04-8.36739924e+00 2.39300602e+00 2.68390216e-02-1.58862068e-05    3
 4.78603122e-09-5.84512948e-13 1.18499465e+04 1.73999551e+01                   4
C3H4-P                  C   3H   4          G    300.00   3500.00 1570.00      1
 6.45797876e+00 1.06371312e-02-3.61161687e-06 5.39412581e-10-2.85851154e-14    2
 1.94136785e+04-1.10770999e+01 1.72714321e+00 2.26902154e-02-1.51273024e-05    3
 5.42930028e-09-8.07229654e-13 2.08991609e+04 1.38804115e+01                   4
C3H4-A                  C   3H   4          G    300.00   3500.00 1420.00      1
 6.37608345e+00 1.10282084e-02-3.89476357e-06 6.16686218e-10-3.59564928e-14    2
 2.00917847e+04-1.13282994e+01 5.08248709e-01 2.75573204e-02-2.13550931e-05    3
 8.81402403e-09-1.47914977e-12 2.17582498e+04 1.90382078e+01                   4
C3H3                    C   3H   3          G    300.00   3500.00  840.00      1
 5.75057757e+00 1.05635748e-02-4.84060955e-06 1.09040069e-09-9.80036131e-14    2
 4.00565408e+04-5.04125036e+00 1.75584160e+00 2.95861270e-02-3.88094528e-05    3
 2.80498001e-08-8.12163438e-12 4.07276565e+04 1.35345457e+01                   4
C3H2                    C   3H   2          G    300.00   3500.00 1260.00      1
 6.42043213e+00 6.05128793e-03-2.30888078e-06 4.10631663e-10-2.84293229e-14    2
 6.08598164e+04-8.32404457e+00 2.15397883e+00 1.95955841e-02-1.84330429e-05    3
 8.94193439e-09-1.72114812e-12 6.19349626e+04 1.32451537e+01                   4
C2H5CHO                 C   3H   6O   1     G    300.00   3500.00 1710.00      1
 9.33264641e+00 1.46861064e-02-4.56011895e-06 5.69517954e-10-1.90907915e-14    2
-2.69164884e+04-2.52385586e+01-9.86882936e-02 3.67477080e-02-2.39124011e-05    3
 8.11426733e-09-1.12212433e-12-2.36909719e+04 2.53220281e+01                   4
CH2CH2CHO               C   3H   5O   1     G    300.00   3500.00  700.00      1
 1.38640407e+00 2.84363937e-02-1.56688639e-05 4.07196319e-09-4.03232081e-13    2
 6.14151621e+02 2.19844215e+01 2.41071813e+00 2.25831705e-02-3.12624277e-06    3
-7.87339030e-09 3.86296559e-12 4.70747652e+02 1.74080454e+01                   4
RALD3                   C   3H   5O   1     G    300.00   3500.00 1140.00      1
-6.08013770e+00 4.60180078e-02-2.61696721e-05 6.65382134e-09-6.35305362e-13    2
-2.14966001e+03 5.90959840e+01 7.04072884e+00-2.01203775e-05 3.44068123e-05    3
-2.87710234e-08 7.13330094e-12-5.14121758e+03-5.92381677e+00                   4
C2H3CHO                 C   3H   4O   1     G    300.00   3500.00 1600.00      1
 9.22597861e+00 1.12038368e-02-3.67974341e-06 5.08180186e-10-2.25803312e-14    2
-1.23719485e+04-2.08137573e+01 8.18907999e-01 3.22215133e-02-2.33838152e-05    3
 8.71821008e-09-1.30539750e-12-9.68168587e+03 2.36968524e+01                   4
CH3COCH3                C   3H   6O   1     G    300.00   3500.00 1790.00      1
 9.79508090e+00 1.35932418e-02-4.01641958e-06 4.43033378e-10-7.94370782e-15    2
-3.07542958e+04-2.70699520e+01-7.54601236e-03 3.54985534e-02-2.23728259e-05    3
 7.27968378e-09-9.62783149e-13-2.72449554e+04 2.59292989e+01                   4
CH3COCH2                C   3H   5O   1     G    300.00   3500.00 1590.00      1
 8.40473974e+00 1.29432016e-02-4.25667165e-06 6.02254308e-10-2.86747777e-14    2
-7.89528966e+03-1.63899873e+01 1.00367425e+00 3.15622343e-02-2.18217968e-05    3
 7.96708666e-09-1.18666729e-12-5.54175084e+03 2.27480013e+01                   4
NC4H10                  C   4H  10          G    300.00   3500.00 1800.00      1
 1.54355394e+01 1.56272489e-02-3.14851571e-06-5.94436194e-11 5.32965842e-14    2
-2.28455274e+04-6.02418014e+01-1.20836791e+00 5.26137097e-02-3.39705664e-05    3
 1.13561307e-08-1.53219985e-12-1.68537208e+04 2.98384973e+01                   4
PC4H9                   C   4H   9          G    300.00   3500.00  950.00      1
 3.94763007e+00 3.16286392e-02-1.12984865e-05 1.11637444e-09 5.54031684e-14    2
 6.05554723e+03 7.76350063e+00-2.76188269e-01 4.94131375e-02-3.93792732e-05    3
 2.08221897e-08-5.13033769e-12 6.85807271e+03 2.79243290e+01                   4
SC4H9                   C   4H   9          G    300.00   3500.00  850.00      1
 3.40122923e+00 3.20901864e-02-1.12255470e-05 9.71712100e-10 8.30726291e-14    2
 4.66283102e+03 1.05291641e+01 2.36336578e-01 4.69837989e-02-3.75083926e-05    3
 2.15857086e-08-5.97986753e-12 5.20086277e+03 2.52835867e+01                   4
IC4H10                  C   4H  10          G    300.00   3500.00 1260.00      1
 5.51955745e+00 3.23747281e-02-1.18655449e-05 1.37455221e-09 1.57072980e-14    2
-1.97025809e+04-6.34483166e+00-1.85965330e+00 5.58007939e-02-3.97537185e-05    3
 1.61301996e-08-2.91200053e-12-1.78430198e+04 3.09610167e+01                   4
IC4H9                   C   4H   9          G    300.00   3500.00 1430.00      1
 7.95880542e+00 2.55088277e-02-8.62221442e-06 8.09648767e-10 4.02033392e-14    2
 3.37759290e+03-1.61084050e+01-1.15582380e+00 5.10042940e-02-3.53657106e-05    3
 1.32774791e-08-2.13948729e-12 5.98437685e+03 3.11244822e+01                   4
TC4H9                   C   4H   9          G    300.00   3500.00 1400.00      1
 7.90871643e+00 2.55264462e-02-8.65284150e-06 8.24420028e-10 3.80550285e-14    2
 8.35470717e+02-1.73299249e+01-1.29900232e+00 5.18342141e-02-3.68397356e-05    3
 1.42467506e-08-2.35878971e-12 3.41363197e+03 3.01901373e+01                   4
IC4H8                   C   4H   8          G    300.00   3500.00 1800.00      1
 7.63433760e+00 2.47722737e-02-1.05415856e-05 2.18152452e-09-1.80119674e-13    2
-6.21385688e+03-1.72949252e+01 7.17301775e-01 4.01434644e-02-2.33509112e-05    3
 6.92571918e-09-8.39035599e-13-3.72372399e+03 2.01415156e+01                   4
IC4H7                   C   4H   7          G    300.00   3500.00  700.00      1
 1.18177126e+00 3.67769034e-02-1.77031335e-05 3.74786261e-09-2.92191278e-13    2
 1.31214242e+04 2.00120535e+01 3.86129974e+00 2.14653122e-02 1.51074192e-05    3
-2.75002829e-08 1.08678607e-11 1.27462902e+04 8.04059820e+00                   4
IC4H7O                  C   4H   7O   1     G    300.00   3500.00 1800.00      1
 1.18822164e+01 1.89918530e-02-7.42296487e-06 1.41442846e-09-1.08683658e-13    2
 1.15971313e+03-3.56333828e+01 1.50010969e+00 4.20632013e-02-2.66490885e-05    3
 8.53521499e-09-1.09768179e-12 4.89727156e+03 2.05567448e+01                   4
C4H8-1                  C   4H   8          G    300.00   3500.00 1800.00      1
 1.03330429e+01 1.99470467e-02-7.40539265e-06 1.30472583e-09-9.09598961e-14    2
-5.56551362e+03-3.07722188e+01-6.91489728e-01 4.44460082e-02-2.78211939e-05    3
 8.86613369e-09-1.14115543e-12-1.59668186e+03 2.88948518e+01                   4
C4H8-2                  C   4H   8          G    300.00   3500.00 1800.00      1
 5.15907751e+00 2.89997624e-02-1.32974550e-05 2.96138882e-09-2.60424337e-13    2
-4.76704818e+03-3.39009988e+00 5.60608160e-01 3.92185832e-02-2.18131390e-05    3
 6.11534585e-09-6.98473924e-13-3.11159921e+03 2.14977755e+01                   4
C4H71-3                 C   4H   7          G    300.00   3500.00 1420.00      1
 8.33017627e+00 1.98466534e-02-6.37614305e-06 5.28653537e-10 3.81102885e-14    2
 1.19533854e+04-1.83767052e+01-1.12550107e+00 4.64823642e-02-3.45124573e-05    3
 1.37381907e-08-2.28751246e-12 1.46387978e+04 3.05571704e+01                   4
C4H71-4                 C   4H   7          G    300.00   3500.00 1530.00      1
 8.45917058e+00 1.93968526e-02-5.99075493e-06 3.82147618e-10 5.73995197e-14    2
 1.98988322e+04-1.80212825e+01-3.29329097e-01 4.23733224e-02-2.85167057e-05    3
 1.01973767e-08-1.54639608e-12 2.25881131e+04 2.81156136e+01                   4
C4H71-O                 C   4H   7O   1     G    300.00   3500.00 1600.00      1
 1.37371780e+01 1.70982840e-02-6.55972505e-06 1.21466080e-09-8.98269511e-14    2
-3.28790330e+01-4.64105988e+01-1.48200932e+00 5.51462524e-02-4.22296954e-05    3
 1.60771484e-08-2.41209064e-12 4.83726092e+03 3.41662559e+01                   4
C4H6                    C   4H   6          G    200.00   3500.00 1800.00      1
 9.30872601e+00 1.50139574e-02-5.06688058e-06 7.84147752e-10-4.70262484e-14    2
 8.60829956e+03-2.47389631e+01 4.65225073e-01 3.46661817e-02-2.14437342e-05    3
 6.84964908e-09-8.89456989e-13 1.17919599e+04 2.31239089e+01                   4
C4H5                    C   4H   5          G    300.00   3500.00 1800.00      1
 1.90192649e+01-1.91794290e-03 4.88814452e-06-1.91833931e-09 2.24139221e-13    2
 3.48592741e+04-7.70423323e+01-2.01742240e-01 4.07954063e-02-3.07063131e-05    3
 1.12647931e-08-1.60685140e-12 4.17788367e+04 2.69857680e+01                   4
C4H4                    C   4H   4          G    300.00   3500.00 1290.00      1
 7.65777095e+00 1.26498264e-02-4.62249002e-06 7.81217249e-10-5.07629295e-14    2
 3.13366017e+04-1.49692649e+01 7.13119750e-01 3.41836286e-02-2.96617949e-05    3
 1.37214265e-08-2.55855542e-12 3.31283217e+04 2.03030642e+01                   4
C4H3                    C   4H   3          G    300.00   3500.00 1590.00      1
 1.30208954e+01 1.53590718e-03 1.80567936e-06-9.30236401e-10 1.18077111e-13    2
 6.01811756e+04-4.25791415e+01 2.34662683e+00 2.83894129e-02-2.35278166e-05    3
 9.69177450e-09-1.55205039e-12 6.35755930e+04 1.38680553e+01                   4
C4H2                    C   4H   2          G    300.00   3500.00  720.00      1
 7.13414721e+00 1.00526312e-02-4.84819237e-06 1.14884615e-09-1.07722848e-13    2
 5.27577825e+04-1.36443509e+01-4.34753587e-01 5.21020801e-02-9.24512109e-05    3
 8.22627522e-08-2.82722735e-11 5.38477042e+04 2.03848055e+01                   4
C6H6                    C   6H   6          G    300.00   3500.00 1410.00      1
 1.15055550e+01 1.99961029e-02-7.07935327e-06 1.10672986e-09-6.24178423e-14    2
 4.11452271e+03-4.24445124e+01-6.99882116e+00 7.24907872e-02-6.29247621e-05    3
 2.75111785e-08-4.74405766e-12 9.33275680e+03 5.31863194e+01                   4
FULVENE                 C   6H   6          G    200.00   3500.00 1560.00      1
 1.44152201e+01 1.47750109e-02-3.90939488e-06 2.82309074e-10 1.62510647e-14    2
 1.91167587e+04-5.54965084e+01-3.67012623e+00 6.11476938e-02-4.84985130e-05    3
 1.93374878e-08-3.03746347e-12 2.47593868e+04 3.97971303e+01                   4
C6H5                    C   6H   5          G    300.00   3500.00 1390.00      1
 1.12331265e+01 1.77269640e-02-6.33615598e-06 1.00236837e-09-5.75481427e-14    2
 3.49856299e+04-3.80075885e+01-6.76261387e+00 6.95132671e-02-6.22206557e-05    3
 2.78054858e-08-4.87825271e-12 3.99884457e+04 5.47375208e+01                   4
C5H6                    C   5H   6          G    200.00   3500.00 1630.00      1
 1.35786775e+01 1.28174233e-02-3.11961760e-06 1.29367868e-10 2.76959074e-14    2
 9.43770546e+03-5.26289111e+01-4.05866650e+00 5.60992491e-02-4.29495186e-05    3
 1.64197159e-08-2.47082373e-12 1.51874796e+04 4.10783322e+01                   4
C5H5                    C   5H   5          G    300.00   3500.00  700.00      1
 4.01652579e+00 2.68451891e-02-1.26423019e-05 2.78092338e-09-2.35299443e-13    2
 2.91110159e+04 1.44025773e+00-2.58737422e+00 6.45817606e-02-9.35063836e-05    3
 7.97943346e-08-2.77400891e-11 3.00355619e+04 3.09448122e+01                   4
MCPTD                   C   6H   8          G    300.00   3500.00 1470.00      1
 1.21408004e+01 2.34281405e-02-7.98703009e-06 1.18908472e-09-6.20202955e-14    2
 7.23040250e+03-4.21606472e+01-5.49894692e+00 7.14274529e-02-5.69659204e-05    3
 2.34017334e-08-3.83968163e-12 1.24164882e+04 4.97368684e+01                   4
C10H8                   C  10H   8          G    300.00   3500.00 1370.00      1
 1.51184866e+01 3.89675471e-02-1.78248571e-05 3.92091997e-09-3.39215370e-13    2
 1.01121550e+04-6.09041302e+01-8.71832459e+00 1.08564076e-01-9.40254364e-05    3
 4.10014938e-08-7.10574345e-12 1.66434413e+04 6.15987891e+01                   4
NC3H7O2                 C   3H   7O   2     G    300.00   3500.00 1650.00      1
 9.25591701e+00 2.27563834e-02-9.54934694e-06 1.92559535e-09-1.53946745e-13    2
-9.34005032e+03-1.86387997e+01 1.92964411e+00 4.05170450e-02-2.56954029e-05    3
 8.44925434e-09-1.14237992e-12-6.92238026e+03 2.03750484e+01                   4
IC3H7O2                 C   3H   7O   2     G    300.00   3500.00 1260.00      1
 7.34738738e+00 2.68252318e-02-1.24179681e-05 2.76645820e-09-2.42147311e-13    2
-1.06484856e+04-8.92587393e+00 1.07341267e+00 4.67426119e-02-3.61291348e-05    3
 1.53120490e-08-2.73135184e-12-9.06744396e+03 2.27924164e+01                   4
C3H7OOH                 C   3H   8O   2     G    300.00   3500.00 1530.00      1
 1.13871490e+01 1.97925486e-02-6.62893833e-06 9.67107057e-10-4.94701006e-14    2
-2.73563036e+04-2.91104764e+01-9.73590419e-01 5.21082072e-02-3.83109566e-05    3
 1.47719080e-08-2.30515654e-12-2.35739173e+04 3.57795698e+01                   4
C3-OQOOH                C   3H   6O   3     G    300.00   3500.00 1350.00      1
 1.12132537e+01 2.34709017e-02-1.13098316e-05 2.59008076e-09-2.30885265e-13    2
-3.91289883e+04-2.66260030e+01 8.46220452e-01 5.41880374e-02-4.54399824e-05    3
 1.94444762e-08-3.35206961e-12-3.63298893e+04 2.65001343e+01                   4
CHOCH2CHO               C   3H   4O   2     G    300.00   3500.00 1370.00      1
 1.06304434e+01 1.18394242e-02-4.21486418e-06 6.67473773e-10-3.88516529e-14    2
-4.37970337e+04-2.83088228e+01-8.46550068e-01 4.53488941e-02-4.09040648e-05    3
 1.85210994e-08-3.29681253e-12-4.06523375e+04 3.06741170e+01                   4
CH2OHCH2CHO             C   3H   6O   2     G    300.00   3500.00 1800.00      1
 1.08721644e+01 1.63593237e-02-6.08637983e-06 1.10130889e-09-8.02911731e-14    2
-4.55272948e+04-2.70748462e+01 2.66105939e+00 3.46062236e-02-2.12921298e-05    3
 6.73306813e-09-8.62479957e-13-4.25712970e+04 1.73653669e+01                   4
CH3CO2H                 C   2H   4O   2     G    300.00   3500.00 1800.00      1
 1.06195335e+01 8.83227209e-03-2.54924796e-06 2.13474537e-10 7.27640500e-15    2
-5.71972748e+04-3.23726626e+01-7.52613302e-01 3.41037094e-02-2.36087790e-05    3
 8.01330086e-09-1.07603281e-12-5.31033019e+04 2.91757681e+01                   4
HCO3                    C   1H   1O   3     G    300.00   3500.00 1490.00      1
 7.67843553e+00 4.62692616e-03-1.54275326e-06 2.12410012e-10-8.98167968e-15    2
-1.61147274e+04-1.27152242e+01 2.31459994e+00 1.90264848e-02-1.60389532e-05    3
 6.69840552e-09-1.09723596e-12-1.45163044e+04 1.53011514e+01                   4
HCO3H                   C   1H   2O   3     G    300.00   3500.00 1750.00      1
 1.00230645e+01 4.43563737e-03-1.56188858e-06 2.43425407e-10-1.38392443e-14    2
-3.81313324e+04-2.33590597e+01 2.47434214e+00 2.16898599e-02-1.63512222e-05    3
 5.87745725e-09-8.18700936e-13-3.54892796e+04 1.72835463e+01                   4
CH2OHCOCH3              C   3H   6O   2     G    300.00   3500.00 1460.00      1
 1.16062108e+01 1.59761338e-02-5.42430613e-06 8.11522207e-10-4.31363898e-14    2
-4.81919049e+04-3.20429601e+01 9.15361391e-01 4.52661321e-02-3.55167701e-05    3
 1.45523733e-08-2.39602186e-12-4.50701769e+04 2.35800151e+01                   4
NC3-QOOH                C   3H   7O   2     G    300.00   3500.00 1800.00      1
 1.29748640e+01 1.76433825e-02-7.16935098e-06 1.42696065e-09-1.14476954e-13    2
-5.86411910e+03-3.67690622e+01 1.55643281e+00 4.30176741e-02-2.83145940e-05    3
 9.25853214e-09-1.20219522e-12-1.75348386e+03 2.50298696e+01                   4
IC3-QOOH                C   3H   7O   2     G    300.00   3500.00 1270.00      1
 1.04498037e+01 2.29490995e-02-1.05757771e-05 2.34172715e-09-2.03669195e-13    2
-5.22299410e+03-2.40008662e+01-1.71110769e-01 5.64007986e-02-5.00856580e-05    3
 2.30818221e-08-4.28636505e-12-2.52528182e+03 2.97774847e+01                   4
NC3-OOQOOH              C   3H   7O   4     G    300.00   3500.00 1260.00      1
 1.11683561e+01 2.95822141e-02-1.42526307e-05 3.27126857e-09-2.92476821e-13    2
-2.00281218e+04-2.06289846e+01 2.57588690e+00 5.68598943e-02-4.67260595e-05    3
 2.04529769e-08-3.70154594e-12-1.78628196e+04 2.28105330e+01                   4
IC3-OOQOOH              C   3H   7O   4     G    300.00   3500.00 1220.00      1
 1.23035626e+01 2.79964881e-02-1.33482909e-05 3.03524082e-09-2.69271163e-13    2
-2.25784830e+04-2.78550806e+01 1.73143834e+00 6.26591905e-02-5.59663676e-05    3
 2.63238073e-08-5.04151840e-12-1.99988847e+04 2.52515835e+01                   4
CH2COOH                 C   2H   3O   2     G    300.00   3500.00 1440.00      1
 1.01170855e+01 5.56298650e-03-8.24127602e-07-2.50445961e-11 1.25384573e-14    2
-3.40138323e+04-2.77197759e+01 4.26277856e-01 3.24818967e-02-2.88646591e-05    3
 1.29566830e-08-2.24123369e-12-3.12228797e+04 2.25664556e+01                   4
IC4-OQOOH               C   4H   8O   3     G    300.00   3500.00 1570.00      1
 1.51567872e+01 2.57227749e-02-1.11020462e-05 2.28943552e-09-1.86269565e-13    2
-4.30658404e+04-4.59844964e+01 9.69279437e-01 6.18692915e-02-4.56369346e-05    3
 1.69539317e-08-2.52138042e-12-3.86109630e+04 2.88616662e+01                   4
NC4-OQOOH               C   4H   8O   3     G    300.00   3500.00 1330.00      1
 1.18153451e+01 3.20093737e-02-1.53334966e-05 3.50316356e-09-3.12136489e-13    2
-4.27660551e+04-2.73083249e+01 2.51946598e+00 5.99669050e-02-4.68645469e-05    3
 1.93082013e-08-3.28300825e-12-4.02933512e+04 2.01899075e+01                   4
C4H9OOH                 C   4H  10O   2     G    300.00   3500.00 1780.00      1
 1.73966955e+01 2.30088682e-02-8.34646818e-06 1.39883156e-09-9.01677199e-14    2
-3.38614044e+04-6.23628989e+01 1.12895114e+00 5.95655972e-02-3.91527005e-05    3
 1.29367463e-08-1.71066136e-12-2.80700874e+04 2.54997631e+01                   4
C5EN-OQOOH-35           C   5H   8O   3     G    300.00   3500.00 1580.00      1
 1.69833158e+01 2.73095006e-02-1.19226835e-05 2.48166871e-09-2.03420335e-13    2
-3.51234524e+04-5.58041843e+01 1.44561311e+00 6.66454568e-02-4.92669457e-05    3
 1.82387414e-08-2.69662803e-12-3.02135384e+04 2.62635808e+01                   4
NC5H10-O                C   5H  10O   1     G    300.00   3500.00 1800.00      1
 1.40073107e+01 3.04405272e-02-1.35854518e-05 2.90305332e-09-2.44985823e-13    2
-2.55455868e+04-5.25239417e+01-3.79263107e+00 6.99959534e-02-4.65483070e-05    3
 1.51115182e-08-1.94060595e-12-1.91376078e+04 4.38130566e+01                   4
NC5-OQOOH               C   5H  10O   3     G    300.00   3500.00 1410.00      1
 1.42172631e+01 3.77707684e-02-1.76257938e-05 3.93443041e-09-3.43954261e-13    2
-4.65061050e+04-3.85369193e+01 2.52749923e+00 7.09332190e-02-5.29049965e-05    3
 2.06149045e-08-3.30148513e-12-4.32095916e+04 2.18759165e+01                   4
NC5H11OOH               C   5H  12O   2     G    300.00   3500.00 1630.00      1
 1.66988185e+01 3.44172714e-02-1.43139763e-05 2.85300857e-09-2.25350885e-13    2
-3.73755763e+04-5.75775300e+01 6.24288977e-02 7.52427673e-02-5.18834510e-05    3
 1.82188469e-08-2.58207456e-12-3.19521133e+04 3.08116404e+01                   4
NC4-QOOH                C   4H   9O   2     G    300.00   3500.00 1760.00      1
 1.83774561e+01 1.83354739e-02-6.23923477e-06 9.66797700e-10-5.61282230e-14    2
-1.29135489e+04-6.55986601e+01 1.19976584e+00 5.73756791e-02-3.95121369e-05    3
 1.35701697e-08-1.84637993e-12-6.86700190e+03 2.69845514e+01                   4
NC4H9-OO                C   4H   9O   2     G    300.00   3500.00 1320.00      1
 8.96630142e+00 3.41074648e-02-1.57640992e-05 3.50715753e-09-3.06662882e-13    2
-1.40847395e+04-1.58347462e+01 9.44281706e-01 5.84166154e-02-4.33881340e-05    3
 1.74586903e-08-2.94899863e-12-1.19669263e+04 2.50940291e+01                   4
IC4H9T-OO               C   4H   9O   2     G    300.00   3500.00 1260.00      1
 9.11667600e+00 3.41757261e-02-1.58797348e-05 3.54686472e-09-3.10976557e-13    2
-1.64591648e+04-1.96564023e+01 4.84069014e-01 6.15808276e-02-4.85048556e-05    3
 2.08088334e-08-3.73597035e-12-1.42837478e+04 2.39860330e+01                   4
IC4T-QOOH               C   4H   9O   2     G    300.00   3500.00 1270.00      1
 1.20890745e+01 3.03954165e-02-1.40883973e-05 3.13822090e-09-2.74437712e-13    2
-1.09705557e+04-3.28537345e+01-4.26302129e-01 6.98139255e-02-6.06456914e-05    3
 2.75777453e-08-5.08536772e-12-7.79165003e+03 3.05171095e+01                   4
IC4P-QOOH               C   4H   9O   2     G    300.00   3500.00 1350.00      1
 1.14809469e+01 3.08095614e-02-1.41939358e-05 3.14755449e-09-2.74422158e-13    2
-7.45268237e+03-2.80879242e+01-1.93281554e-01 6.53998681e-02-5.26276099e-05    3
 2.21271466e-08-3.78916144e-12-4.30064068e+03 3.17369695e+01                   4
IC4H9P-OO               C   4H   9O   2     G    300.00   3500.00 1380.00      1
 8.54295878e+00 3.45220761e-02-1.59311934e-05 3.53852644e-09-3.08950026e-13    2
-1.29532174e+04-1.39825096e+01 7.00555087e-01 5.72536810e-02-4.06394596e-05    3
 1.54748869e-08-2.47133417e-12-1.07887140e+04 2.63784637e+01                   4
NC4-OOQOOH              C   4H   9O   4     G    300.00   3500.00 1230.00      1
 1.51474115e+01 3.37812806e-02-1.58996821e-05 3.57608780e-09-3.14486500e-13    2
-2.85698877e+04-4.24732212e+01 1.10123473e+00 7.94599042e-02-7.16053206e-05    3
 3.37688458e-08-6.45122593e-12-2.51145282e+04 2.81992198e+01                   4
IC4T-OOQOOH             C   4H   9O   4     G    300.00   3500.00 1240.00      1
 1.39939781e+01 3.54845225e-02-1.68915062e-05 3.83671085e-09-3.40131623e-13    2
-2.83614519e+04-3.70531084e+01 1.55094394e+00 7.56233423e-02-6.54465301e-05    3
 2.99415625e-08-5.60320654e-12-2.52755794e+04 2.56539769e+01                   4
IC4P-OOQOOH             C   4H   9O   4     G    300.00   3500.00 1290.00      1
 1.30518456e+01 3.65484776e-02-1.74274761e-05 3.96741885e-09-3.52551959e-13    2
-2.47096142e+04-3.04334752e+01 1.64511772e+00 7.19181763e-02-5.85550328e-05    3
 2.52219701e-08-4.47165103e-12-2.17666784e+04 2.75020274e+01                   4
C5EN-QOOH               C   5H   9O   2     G    300.00   3500.00 1420.00      1
 1.28791282e+01 3.32930438e-02-1.55378912e-05 3.46674357e-09-3.02869760e-13    2
 3.23011696e+03-3.38507217e+01 1.34404403e+00 6.57862385e-02-4.98616884e-05    3
 1.95812024e-08-3.13992237e-12 6.50608086e+03 2.58442478e+01                   4
C5EN-OO                 C   5H   9O   2     G    300.00   3500.00 1280.00      1
 1.00840313e+01 3.69913058e-02-1.74216198e-05 3.93130809e-09-3.47257470e-13    2
-8.98414916e+02-1.96513594e+01 4.09897394e-01 6.72229742e-02-5.28493562e-05    3
 2.23832541e-08-3.95115317e-12 1.57816335e+03 2.94089017e+01                   4
C5EN-OOQOOH-35          C   5H   9O   4     G    300.00   3500.00 1160.00      1
 1.36699768e+01 4.21231927e-02-2.15503705e-05 5.21806313e-09-4.87292988e-13    2
-1.42354804e+04-3.35883377e+01 5.24578548e-01 8.74521521e-02-8.01654042e-05    3
 3.89048641e-08-7.74737940e-12-1.11857480e+04 3.17816499e+01                   4
NC5H12OO                C   5H  11O   2     G    300.00   3500.00 1300.00      1
 1.06544843e+01 4.16170567e-02-1.93382878e-05 4.32113973e-09-3.79088258e-13    2
-1.98652038e+04-2.50234562e+01 3.19664945e-01 7.34165010e-02-5.60299543e-05    3
 2.31373790e-08-3.99759580e-12-1.71781508e+04 2.75475606e+01                   4
NC5-QOOH                C   5H  11O   2     G    300.00   3500.00 1300.00      1
 1.36538185e+01 3.77860044e-02-1.75151101e-05 3.90394490e-09-3.41708634e-13    2
-1.43879857e+04-3.94678771e+01-5.74282925e-01 8.15647781e-02-6.80290797e-05    3
 2.98085447e-08-5.32336244e-12-1.06886793e+04 3.29074330e+01                   4
NC5-OOQOOH              C   5H  11O   4     G    300.00   3500.00 1270.00      1
 1.54638471e+01 4.30531989e-02-2.04284739e-05 4.63174757e-09-4.10272033e-13    2
-3.17413364e+04-4.31406891e+01 1.43265575e+00 8.72459276e-02-7.26246102e-05    3
 3.20312942e-08-5.80388357e-12-2.81774138e+04 2.79053903e+01                   4
C4H6O2                  C   4H   6O   2     G    300.00   3500.00 1800.00      1
 7.01919732e+00 2.89919931e-02-1.39811142e-05 3.22750413e-09-2.90888748e-13    2
-4.36055716e+04-7.47847768e+00 9.15158131e-01 4.25565247e-02-2.52848905e-05    3
 7.41408794e-09-8.72358721e-13-4.14081175e+04 2.55578558e+01                   4
C4H8O                   C   4H   8O   1     G    300.00   3500.00 1800.00      1
 1.12815969e+01 2.48463755e-02-1.13234737e-05 2.47070049e-09-2.12413611e-13    2
-2.03756677e+04-3.84267219e+01-2.94845096e+00 5.64687040e-02-3.76754141e-05    3
 1.22306784e-08-1.56796610e-12-1.52528505e+04 3.85892654e+01                   4
C5H8O                   C   5H   8O   1     G    300.00   3500.00 1330.00      1
 6.70800638e+00 3.65243787e-02-1.77765832e-05 4.15639182e-09-3.79163349e-13    2
-5.52771767e+03-9.67918152e+00-5.12640157e+00 7.21165831e-02-5.79181670e-05    3
 2.42774865e-08-4.16132400e-12-2.37976515e+03 5.07899198e+01                   4
RNC3OHOOX               C   3H   7O   3     G    300.00   3500.00 1800.00      1
 3.74667467e+01 1.57251514e-02-1.09732354e-05 3.61008676e-09-4.15087623e-13    2
-5.05275841e+04-1.70384642e+02-4.06427157e+00 1.08016303e-01-8.78825284e-05    3
 3.20950101e-08-4.37132697e-12-3.55764175e+04 5.43898919e+01                   4
QNC3OHOOX               C   3H   7O   3     G    300.00   3500.00 1800.00      1
 3.65507341e+01 1.64042496e-02-1.14786834e-05 3.72939233e-09-4.24701786e-13    2
-4.45414868e+04-1.61156405e+02-1.59743962e+00 1.01177969e-01-8.21234495e-05    3
 2.98941205e-08-4.05869181e-12-3.08081442e+04 4.53094695e+01                   4
ZNC3OHOOX               C   3H   7O   5     G    300.00   3500.00 1140.00      1
 2.54947967e+01 2.87030621e-02-3.65256446e-06-1.12208373e-09 2.39300330e-13    2
-5.46882914e+04-8.79716172e+01-1.83124933e+00 1.24583925e-01-1.29811595e-04    3
 7.26551271e-08-1.59399126e-11-4.84579529e+04 4.74412433e+01                   4
KEHYNC3OH               C   3H   6O   4     G    300.00   3500.00  990.00      1
 2.03864539e+01 2.59482566e-02 2.17638899e-06-3.94711697e-09 6.27440524e-13    2
-7.09480078e+04-6.09332078e+01-1.73111502e+00 1.15312171e-01-1.33223482e-04    3
 8.72312472e-08-2.23973989e-11-6.65687292e+04 4.55489880e+01                   4
C3OHCYETH               C   3H   6O   2     G    200.00   3500.00 1670.00      1
 1.35374615e+01 1.18925377e-02-2.94432386e-06 1.64021062e-10 1.84650891e-14    2
-3.51827728e+04-4.61976510e+01-8.63498967e-01 4.63858562e-02-3.39263465e-05    3
 1.25320940e-08-1.83304283e-12-3.03728520e+04 3.06638116e+01                   4
RBU1OOX                 C   4H   9O   3     G    300.00   3500.00 1670.00      1
 1.45390313e+01 2.69797342e-02-1.09312492e-05 2.12602312e-09-1.64284691e-13    2
-3.56893367e+04-4.22613598e+01 3.26237582e+00 5.39896876e-02-3.51916863e-05    3
 1.18108284e-08-1.61410584e-12-3.19229337e+04 1.79249199e+01                   4
QBU1OOX                 C   4H   9O   3     G    300.00   3500.00 1270.00      1
 9.44680429e+00 1.40890834e-02-6.70668655e-06 1.51288708e-09-1.32818601e-13    2
 1.91332918e+04-2.81812909e+01-5.88861866e+00 6.23896281e-02-6.37545740e-05    3
 3.14592847e-08-6.02777876e-12 2.30284892e+04 4.94686853e+01                   4
ZBU1OOX                 C   4H   9O   5     G    300.00   3500.00 1410.00      1
 1.71509970e+01 3.21642998e-02-1.45265252e-05 3.16055989e-09-2.71089898e-13    2
-4.87167966e+04-4.94521673e+01 4.90929019e+00 6.68925459e-02-5.14714679e-05    3
 2.06286179e-08-3.36826331e-12-4.52646353e+04 1.38131159e+01                   4
KEHYBU1                 C   4H   8O   4     G    300.00   3500.00 1200.00      1
 1.50812006e+01 2.99746625e-02-1.37944077e-05 3.03171339e-09-2.60935165e-13    2
-6.34178096e+04-4.27051085e+01-4.53521769e+00 9.53627234e-02-9.55294838e-05    3
 4.84400890e-08-9.72101341e-12-5.87098692e+04 5.55092662e+01                   4
C4OHCYETH               C   4H   8O   2     G    300.00   3500.00 1740.00      1
 1.55057880e+01 1.98739170e-02-6.85214241e-06 1.07267976e-09-6.29459251e-14    2
-5.34275304e+04-5.89096443e+01-4.24192759e+00 6.52709644e-02-4.59875281e-05    3
 1.60670804e-08-2.21731383e-12-4.65553254e+04 4.72996339e+01                   4
RPENT1OOX               C   5H  11O   3     G    300.00   3500.00 1690.00      1
 2.06735989e+01 3.07534954e-02-1.19967931e-05 2.22747833e-09-1.63728718e-13    2
-5.79272417e+04-7.43003333e+01 2.17872322e+00 7.45283490e-02-5.08502135e-05    3
 1.75542714e-08-2.43100580e-12-5.16759738e+04 2.46315395e+01                   4
QPENT1OOX               C   5H  11O   3     G    300.00   3500.00 1590.00      1
 1.99691796e+01 3.07316175e-02-1.29590636e-05 2.61520597e-09-2.08804239e-13    2
-3.62027685e+04-6.96874712e+01 1.91284963e+00 7.61563469e-02-5.58125819e-05    3
 2.05831382e-08-3.03395081e-12-3.04608556e+04 2.57972176e+01                   4
ZPENT1OOX               C   5H  11O   5     G    300.00   3500.00 1380.00      1
 2.07046201e+01 3.73731215e-02-1.71331760e-05 3.77821831e-09-3.27723703e-13    2
-5.43479695e+04-6.52594396e+01 3.53770720e+00 8.71322893e-02-7.12192280e-05    3
 2.99067458e-08-5.06115260e-12-4.96099015e+04 2.30901711e+01                   4
KEHYP1OH                C   5H  10O   4     G    300.00   3500.00 1560.00      1
 1.98034559e+01 3.06181813e-02-1.26872565e-05 2.52829397e-09-2.00061856e-13    2
-6.77003658e+04-6.61563442e+01 2.43438013e+00 7.51542730e-02-5.55104216e-05    3
 2.08287919e-08-3.13283395e-12-6.22812142e+04 2.53631878e+01                   4
C5OHCYETH               C   5H  10O   2     G    300.00   3500.00 1760.00      1
 1.88847141e+01 2.52072174e-02-8.75962755e-06 1.38787272e-09-8.30557860e-14    2
-5.99419471e+04-8.09815610e+01-5.15784759e+00 7.98494032e-02-5.53296722e-05    3
 1.90280412e-08-2.58876153e-12-5.14789654e+04 4.86014936e+01                   4
RC6OHOOX                C   6H  13O   3     G    300.00   3500.00 1800.00      1
 3.74667467e+01 1.57251514e-02-1.09732354e-05 3.61008676e-09-4.15087623e-13    2
-5.05275841e+04-1.70384642e+02-4.06427157e+00 1.08016303e-01-8.78825284e-05    3
 3.20950101e-08-4.37132697e-12-3.55764175e+04 5.43898919e+01                   4
QC6OHOOX                C   6H  13O   3     G    300.00   3500.00 1800.00      1
 3.65507341e+01 1.64042496e-02-1.14786834e-05 3.72939233e-09-4.24701786e-13    2
-4.45414868e+04-1.61156405e+02-1.59743962e+00 1.01177969e-01-8.21234495e-05    3
 2.98941205e-08-4.05869181e-12-3.08081442e+04 4.53094695e+01                   4
ZC6OHOOX                C   6H  13O   5     G    300.00   3500.00 1140.00      1
 2.54947967e+01 2.87030621e-02-3.65256446e-06-1.12208373e-09 2.39300330e-13    2
-5.46882914e+04-8.79716172e+01-1.83124933e+00 1.24583925e-01-1.29811595e-04    3
 7.26551271e-08-1.59399126e-11-4.84579529e+04 4.74412433e+01                   4
KEHYC6OH                C   6H  12O   4     G    300.00   3500.00  990.00      1
 2.03864539e+01 2.59482566e-02 2.17638899e-06-3.94711697e-09 6.27440524e-13    2
-7.09480078e+04-6.09332078e+01-1.73111502e+00 1.15312171e-01-1.33223482e-04    3
 8.72312472e-08-2.23973989e-11-6.65687292e+04 4.55489880e+01                   4
C6OHCYETH               C   6H  12O   2     G    300.00   3500.00 1760.00      1
 1.88847141e+01 2.52072174e-02-8.75962755e-06 1.38787272e-09-8.30557860e-14    2
-5.99419471e+04-8.09815610e+01-5.15784759e+00 7.98494032e-02-5.53296722e-05    3
 1.90280412e-08-2.58876153e-12-5.14789654e+04 4.86014936e+01                   4
RALD3OO                 C   3H   5O   3     G    300.00   3500.00 1800.00      1
 1.58771652e+01 1.28699625e-02-5.29703455e-06 1.04001972e-09-8.12487350e-14    2
-2.38887628e+04-5.44666560e+01 3.38301201e+00 4.06347474e-02-2.84343553e-05    3
 9.60939777e-09-1.27144013e-12-1.93908676e+04 1.31543075e+01                   4
QALD3OO                 C   3H   5O   3     G    300.00   3500.00 1300.00      1
 1.09154406e+01 2.11069280e-02-1.04347914e-05 2.43633202e-09-2.20224994e-13    2
-1.35446351e+04-2.42468422e+01 1.81101369e+00 4.91205491e-02-4.27582004e-05    3
 1.90124392e-08-3.40793791e-12-1.11774841e+04 2.20654309e+01                   4
ZALD3OO                 C   3H   5O   5     G    300.00   3500.00 1800.00      1
 2.14549181e+01 1.08256429e-02-3.75393411e-06 5.88014390e-10-3.47283349e-14    2
-3.59900206e+04-7.93559827e+01 5.41191672e+00 4.64767571e-02-3.34631960e-05    3
 1.15914447e-08-1.56298255e-12-3.02145401e+04 7.47208774e+00                   4
ETC3H4O2                C   3H   4O   2     G    300.00   3500.00 1240.00      1
 1.02920433e+01 1.38871288e-02-6.12561891e-06 1.30548810e-09-1.09965724e-13    2
-3.57026990e+04-2.69350056e+01 1.17378026e-01 4.67086296e-02-4.58290473e-05    3
 2.26514173e-08-4.41358049e-12-3.31793820e+04 2.43405590e+01                   4
KEA3B3L                 C   3H   4O   4     G    300.00   3500.00 1500.00      1
 1.56495509e+01 1.47904687e-02-6.84032207e-06 1.49167075e-09-1.26830295e-13    2
-4.74213142e+04-4.92482800e+01 1.41905654e+00 5.27384538e-02-4.47883071e-05    3
 1.83574419e-08-2.93779215e-12-4.31521659e+04 2.51755985e+01                   4
RALD4OOX                C   4H   7O   3     G    300.00   3500.00 1060.00      1
 1.47280764e+01 1.68541720e-02-7.08657288e-07-1.32138230e-09 2.25378312e-13    2
-2.49490049e+04-4.17540778e+01-2.51677560e+00 8.19290854e-02-9.27957989e-05    3
 5.65950589e-08-1.34341597e-11-2.12930963e+04 4.24472036e+01                   4
QA4X                    C   4H   7O   3     G    300.00   3500.00 1020.00      1
 1.57879646e+01 1.38870675e-02 1.11593595e-06-1.77746718e-09 2.67503325e-13    2
-1.92489294e+04-4.33532544e+01-6.30635463e-01 7.82737344e-02-9.35703389e-05    3
 6.01089870e-08-1.49007452e-11-1.58995350e+04 3.61821315e+01                   4
ZA4X                    C   4H   7O   5     G    300.00   3500.00 1030.00      1
 2.21686908e+01 9.17757366e-03 7.13282519e-06-4.12053823e-09 5.56292343e-13    2
-3.97162882e+04-7.35383795e+01-2.33834089e+00 1.04350512e-01-1.31468542e-04    3
 8.55890844e-08-2.12178879e-11-3.46678396e+04 4.54182805e+01                   4
KEA4X                   C   4H   6O   4     G    300.00   3500.00  980.00      1
 1.51486381e+01 1.43075631e-02 4.47525116e-07-1.46947381e-09 2.26509050e-13    2
-1.74087245e+04-3.88103570e+01 7.77077995e-01 7.29669921e-02-8.93373151e-05    3
 5.96086488e-08-1.53546447e-11-1.45918987e+04 3.02337685e+01                   4
ETALD4X                 C   4H   6O   2     G    300.00   3500.00 1200.00      1
 9.47104175e+00 1.56985812e-02-7.47624864e-06 1.72107270e-09-1.55288678e-13    2
-3.54471815e+04-2.25395264e+01 7.88831220e-02 4.70057766e-02-4.66102429e-05    3
 2.34621806e-08-4.68468617e-12-3.31930634e+04 2.44846028e+01                   4
CH3COCHO                C   3H   4O   2     G    300.00   3500.00 1370.00      1
 1.06304434e+01 1.18394242e-02-4.21486418e-06 6.67473773e-10-3.88516529e-14    2
-4.37970337e+04-2.83088228e+01-8.46550068e-01 4.53488941e-02-4.09040648e-05    3
 1.85210994e-08-3.29681253e-12-4.06523375e+04 3.06741170e+01                   4
RALD5XOO                C   5H   9O   3     G    300.00   3500.00 1240.00      1
 5.00092597e+01-5.34134319e-02 6.46290192e-05-2.28767019e-08 2.64030379e-12    2
-4.06673535e+04-2.20829578e+02-1.12640291e+01 1.44242338e-01-1.74470703e-04    3
 1.05671536e-07-2.32766796e-11-2.54715779e+04 8.79592024e+01                   4
QA5X                    C   5H   9O   3     G    300.00   3500.00 1020.00      1
 3.16179270e+01-1.36493871e-02 3.39152641e-05-1.31900624e-08 1.56959108e-12    2
-3.26152699e+04-1.14322462e+02-3.56697921e+00 1.24330637e-01-1.68996536e-04    3
 1.19432029e-07-3.09358236e-11-2.54375491e+04 5.61211251e+01                   4
ZA5X                    C   5H   9O   5     G    300.00   3500.00 1030.00      1
 4.82844916e+01-4.15707461e-02 6.14657160e-05-2.30375139e-08 2.73823900e-12    2
-5.69207575e+04-1.98450742e+02-1.56034012e+01 2.06537576e-01-2.99857083e-04    3
 2.10828375e-07-5.40253263e-11-4.37598516e+04 1.11659860e+02                   4
KEA5X                   C   5H   8O   4     G    300.00   3500.00  890.00      1
 2.81159854e+01-1.51101034e-02 3.53666263e-05-1.35086152e-08 1.59169636e-12    2
 3.74972700e+04-9.42664383e+01 2.11579827e-01 1.10302955e-01-1.76003697e-04    3
 1.44821215e-07-4.28829751e-11 4.24642542e+04 3.71043815e+01                   4
RALD6XOO                C   6H  11O   3     G    300.00   3500.00 1240.00      1
 5.00092597e+01-5.34134319e-02 6.46290192e-05-2.28767019e-08 2.64030379e-12    2
-4.06673535e+04-2.20829578e+02-1.12640291e+01 1.44242338e-01-1.74470703e-04    3
 1.05671536e-07-2.32766796e-11-2.54715779e+04 8.79592024e+01                   4
QA6X                    C   6H  11O   3     G    300.00   3500.00 1020.00      1
 3.16179270e+01-1.36493871e-02 3.39152641e-05-1.31900624e-08 1.56959108e-12    2
-3.26152699e+04-1.14322462e+02-3.56697921e+00 1.24330637e-01-1.68996536e-04    3
 1.19432029e-07-3.09358236e-11-2.54375491e+04 5.61211251e+01                   4
ZA6X                    C   6H  11O   5     G    300.00   3500.00 1030.00      1
 4.82844916e+01-4.15707461e-02 6.14657160e-05-2.30375139e-08 2.73823900e-12    2
-5.69207575e+04-1.98450742e+02-1.56034012e+01 2.06537576e-01-2.99857083e-04    3
 2.10828375e-07-5.40253263e-11-4.37598516e+04 1.11659860e+02                   4
KEA6X                   C   6H  10O   4     G    300.00   3500.00  890.00      1
 2.81159854e+01-1.51101034e-02 3.53666263e-05-1.35086152e-08 1.59169636e-12    2
 3.74972700e+04-9.42664383e+01 2.11579827e-01 1.10302955e-01-1.76003697e-04    3
 1.44821215e-07-4.28829751e-11 4.24642542e+04 3.71043815e+01                   4
ETALD6X                 C   6H  10O   2     G    300.00   3500.00 1200.00      1
 9.47104175e+00 1.56985812e-02-7.47624864e-06 1.72107270e-09-1.55288678e-13    2
-3.54471815e+04-2.25395264e+01 7.88831220e-02 4.70057766e-02-4.66102429e-05    3
 2.34621806e-08-4.68468617e-12-3.31930634e+04 2.44846028e+01                   4
RIBALDGOO               C   4H   7O   3     G    300.00   3500.00 1090.00      1
 1.33433410e+01 1.84987684e-02-1.85145411e-06-9.50436871e-10 1.82631111e-13    2
-2.33799979e+04-3.43356019e+01-3.50808847e+00 8.03388765e-02-8.69525203e-05    3
 5.10991449e-08-1.17553464e-11-1.97063863e+04 4.84150215e+01                   4
RIBALDBOO               C   4H   7O   3     G    300.00   3500.00 1060.00      1
 1.47280764e+01 1.68541720e-02-7.08657288e-07-1.32138230e-09 2.25378312e-13    2
-2.49490049e+04-4.17540778e+01-2.51677560e+00 8.19290854e-02-9.27957989e-05    3
 5.65950589e-08-1.34341597e-11-2.12930963e+04 4.24472036e+01                   4
QIBALDG2                C   4H   7O   3     G    300.00   3500.00  980.00      1
 1.67965092e+01 1.08043145e-02 4.76342236e-06-3.20053212e-09 4.44231176e-13    2
-2.25755349e+04-5.02646438e+01-3.01325452e-01 8.05913947e-02-1.02053537e-04    3
 6.94640662e-08-1.80926561e-11-1.92243593e+04 3.18771024e+01                   4
QIBALDG3                C   4H   7O   3     G    300.00   3500.00 1050.00      1
 1.47854636e+01 1.55385627e-02-2.73488914e-07-1.29944011e-09 2.11492588e-13    2
-1.68282753e+04-3.82904654e+01-2.35309170e+00 8.08282972e-02-9.35445382e-05    3
 5.79202737e-08-1.38884393e-11-1.32291787e+04 4.52293499e+01                   4
QIBALDB3                C   4H   7O   3     G    300.00   3500.00 1020.00      1
 1.57879646e+01 1.38870675e-02 1.11593595e-06-1.77746718e-09 2.67503325e-13    2
-1.92489294e+04-4.33532544e+01-6.30635463e-01 7.82737344e-02-9.35703389e-05    3
 6.01089870e-08-1.49007452e-11-1.58995350e+04 3.61821315e+01                   4
ETIBALDGB               C   4H   6O   2     G    300.00   3500.00 1200.00      1
 9.47104175e+00 1.56985812e-02-7.47624864e-06 1.72107270e-09-1.55288678e-13    2
-3.54471815e+04-2.25395264e+01 7.88831220e-02 4.70057766e-02-4.66102429e-05    3
 2.34621806e-08-4.68468617e-12-3.31930634e+04 2.44846028e+01                   4
ETIBALDGG               C   4H   6O   2     G    300.00   3500.00 1200.00      1
 9.47104175e+00 1.56985812e-02-7.47624864e-06 1.72107270e-09-1.55288678e-13    2
-3.54471815e+04-2.25395264e+01 7.88831220e-02 4.70057766e-02-4.66102429e-05    3
 2.34621806e-08-4.68468617e-12-3.31930634e+04 2.44846028e+01                   4
ZIBALDG2                C   4H   7O   5     G    300.00   3500.00 1030.00      1
 2.21686908e+01 9.17757366e-03 7.13282519e-06-4.12053823e-09 5.56292343e-13    2
-3.97162882e+04-7.35383795e+01-2.33834089e+00 1.04350512e-01-1.31468542e-04    3
 8.55890844e-08-2.12178879e-11-3.46678396e+04 4.54182805e+01                   4
ZIBALDG3                C   4H   7O   5     G    300.00   3500.00 1080.00      1
 1.90668847e+01 1.53920270e-02 1.15889307e-06-1.93814966e-09 2.92451704e-13    2
-3.52242061e+04-5.68408622e+01-2.45362858e+00 9.50976317e-02-1.09543336e-04    3
 6.63965594e-08-1.55257680e-11-3.05757753e+04 4.86394153e+01                   4
ZIBALDB3                C   4H   7O   5     G    300.00   3500.00 1080.00      1
 1.90668847e+01 1.53920270e-02 1.15889307e-06-1.93814966e-09 2.92451704e-13    2
-3.52242061e+04-5.68408622e+01-2.45362858e+00 9.50976317e-02-1.09543336e-04    3
 6.63965594e-08-1.55257680e-11-3.05757753e+04 4.86394153e+01                   4
KIA4G2                  C   4H   6O   4     G    300.00   3500.00 1800.00      1
 2.35089834e+01 2.55786937e-03-1.96914986e-06 1.09436504e-09-1.65130016e-13    2
-5.44782537e+04-9.88855006e+01-1.84484574e+00 5.88997119e-02-4.89206853e-05    3
 1.84838226e-08-2.58033246e-12-4.53508752e+04 3.83347117e+01                   4
NEOC5H10-O              C   5H  10O   1     G    300.00   3500.00 1470.00      1
 1.29296113e+01 3.16150586e-02-1.35584955e-05 2.81753122e-09-2.32686212e-13    2
-2.37933927e+04-4.88968600e+01-6.91462643e+00 8.56129843e-02-6.86584196e-05    3
 2.78061590e-08-4.48245283e-12-1.79591868e+04 5.44853544e+01                   4
NEOC5-OQOOH             C   5H  10O   3     G    300.00   3500.00 1690.00      1
 2.24459975e+01 2.37621197e-02-8.83880918e-06 1.53829914e-09-1.04514649e-13    2
-5.03880263e+04-8.77405842e+01 1.27283517e+00 7.38761133e-02-5.33186852e-05    3
 1.90846013e-08-2.70012148e-12-4.32314975e+04 2.55178470e+01                   4
NEOC5H11-OO             C   5H  11O   2     G    300.00   3500.00 1660.00      1
 1.69989725e+01 3.01601512e-02-1.19254906e-05 2.25822396e-09-1.69878978e-13    2
-2.10464566e+04-6.14617694e+01 1.07910956e+00 6.85212668e-02-4.65891492e-05    3
 1.61793720e-08-2.26643742e-12-1.57610621e+04 2.34108335e+01                   4
NEOC5-QOOH              C   5H  11O   2     G    300.00   3500.00 1630.00      1
 1.86197572e+01 2.85111334e-02-1.13969269e-05 2.18137062e-09-1.65768739e-13    2
-1.50391461e+04-6.74883963e+01 1.48070264e+00 7.05701629e-02-5.01015553e-05    3
 1.80114845e-08-2.59370031e-12-9.45181433e+03 2.35714339e+01                   4
NEOC5-OOQOOH            C   5H  11O   4     G    300.00   3500.00 1800.00      1
 2.53088265e+01 2.46008498e-02-8.38585078e-06 1.28446276e-09-7.25492644e-14    2
-3.52662106e+04-9.88693070e+01 2.93992997e+00 7.43095087e-02-4.98097332e-05    3
 1.66266415e-08-2.20340742e-12-2.72134078e+04 2.21958274e+01                   4
CYC6-OO                 C   6H  11O   2     G    300.00   3500.00 1800.00      1
 1.87814636e+01 3.54361897e-02-1.49718764e-05 3.04328229e-09-2.46478261e-13    2
-1.95252836e+04-7.87240961e+01-6.50623583e+00 9.16310773e-02-6.18009494e-05    3
 2.03873834e-08-2.65538120e-12-1.04217118e+04 5.81382086e+01                   4
CYC6-QOOH-2             C   6H  11O   2     G    300.00   3500.00 1800.00      1
 1.91384114e+01 3.64873128e-02-1.63613005e-05 3.53264682e-09-3.02111809e-13    2
-1.43294339e+04-7.86383458e+01-4.87015373e+00 8.98396797e-02-6.08216063e-05    3
 1.99994267e-08-2.58916458e-12-5.68635041e+03 5.13010171e+01                   4
CYC6-QOOH-3             C   6H  11O   2     G    300.00   3500.00 1800.00      1
 2.09300716e+01 3.28719806e-02-1.40160786e-05 2.89193659e-09-2.38539859e-13    2
-1.52994540e+04-8.89349599e+01-7.04914209e+00 9.50480110e-02-6.58294373e-05    3
 2.20820695e-08-2.90383609e-12-5.22693705e+03 6.24943814e+01                   4
CYC6-QOOH-4             C   6H  11O   2     G    300.00   3500.00 1800.00      1
 2.09300716e+01 3.28719806e-02-1.40160786e-05 2.89193659e-09-2.38539859e-13    2
-1.52994540e+04-8.89349599e+01-7.04914209e+00 9.50480110e-02-6.58294373e-05    3
 2.20820695e-08-2.90383609e-12-5.22693705e+03 6.24943814e+01                   4
CYC6H10-O-12            C   6H  10O   1     G    300.00   3500.00 1800.00      1
 2.29323137e+01 2.20056630e-02-7.35242861e-06 1.07816550e-09-5.64637362e-14    2
-2.79806185e+04-1.10525182e+02-1.05629253e+01 9.64395276e-02-6.93806491e-05    3
 2.40515805e-08-3.24721582e-12-1.59223324e+04 7.07580390e+01                   4
CYC6H10-O-13            C   6H  10O   1     G    300.00   3500.00 1800.00      1
 2.18028749e+01 2.41377149e-02-8.73116363e-06 1.46035059e-09-9.51861242e-14    2
-2.87387506e+04-1.06217600e+02-1.25990105e+01 1.00586349e-01-7.24383588e-05    3
 2.50556081e-08-3.37230522e-12-1.63540718e+04 7.99725804e+01                   4
CYC6H10-O-14            C   6H  10O   1     G    300.00   3500.00 1800.00      1
 2.14079716e+01 2.50825212e-02-9.38037933e-06 1.64524949e-09-1.14247149e-13    2
-3.89741865e+04-1.05728301e+02-1.45960527e+01 1.05091464e-01-7.60544985e-05    3
 2.63393677e-08-3.54398579e-12-2.60127377e+04 8.91329893e+01                   4
CYC6H10-ONE             C   6H  10O   1     G    300.00   3500.00 1800.00      1
 1.15965456e+01 4.02887877e-02-1.86685801e-05 4.15568325e-09-3.64030600e-13    2
-3.62221504e+04-4.27468590e+01-6.46490405e+00 8.04253425e-02-5.21157091e-05    3
 1.65435088e-08-2.08456193e-12-2.97200285e+04 5.50054745e+01                   4
C5H9CHO                 C   6H  10O   1     G    300.00   3500.00 1100.00      1
 9.07727149e+00 2.66919106e-02-7.89644734e-06 7.31227443e-10 1.61730797e-14    2
-1.68606426e+04-1.54909484e+01-3.32869078e-01 6.09106036e-02-5.45583014e-05    3
 2.90111390e-08-6.41107955e-12-1.47904117e+04 3.08044225e+01                   4
CYC6-OOQOOH-2           C   6H  11O   4     G    300.00   3500.00 1770.00      1
 2.93742106e+01 2.67859027e-02-9.56347572e-06 1.54086137e-09-9.31288498e-14    2
-3.55499006e+04-1.29752722e+02-4.99061868e+00 1.04446534e-01-7.53775698e-05    3
 2.63295974e-08-3.59436275e-12-2.33847511e+04 5.56593291e+01                   4
CYC6-OOQOOH-3           C   6H  11O   4     G    300.00   3500.00 1770.00      1
 2.93742106e+01 2.67859027e-02-9.56347572e-06 1.54086137e-09-9.31288498e-14    2
-3.55499006e+04-1.29752722e+02-4.99061868e+00 1.04446534e-01-7.53775698e-05    3
 2.63295974e-08-3.59436275e-12-2.33847511e+04 5.56593291e+01                   4
CYC6-OOQOOH-4           C   6H  11O   4     G    300.00   3500.00 1770.00      1
 2.93742106e+01 2.67859027e-02-9.56347572e-06 1.54086137e-09-9.31288498e-14    2
-3.55499006e+04-1.30447236e+02-4.99061868e+00 1.04446534e-01-7.53775698e-05    3
 2.63295974e-08-3.59436275e-12-2.33847511e+04 5.49648151e+01                   4
CYC6-OQOOH-2            C   6H  10O   3     G    300.00   3500.00 1460.00      1
 1.17655252e+01 3.67451381e-02-1.42717430e-05 2.74140392e-09-2.13135444e-13    2
-3.59903396e+04-5.10812548e+01-1.06696445e+01 9.82113564e-02-7.74219672e-05    3
 3.15771228e-08-5.15075853e-12-2.94392700e+04 6.56457557e+01                   4
CYC6-OQOOH-3            C   6H  10O   3     G    300.00   3500.00 1460.00      1
 1.16022426e+01 3.57303644e-02-1.34415869e-05 2.50437418e-09-1.89510245e-13    2
-3.63821559e+04-4.91587855e+01-8.02402170e+00 8.95009515e-02-6.86853407e-05    3
 2.77298326e-08-4.50893805e-12-3.06512867e+04 5.29538882e+01                   4
CYC6-OQOOH-4            C   6H  10O   3     G    300.00   3500.00 1460.00      1
 1.16022426e+01 3.57303644e-02-1.34415869e-05 2.50437418e-09-1.89510245e-13    2
-3.63821559e+04-4.98532999e+01-8.02402170e+00 8.95009515e-02-6.86853407e-05    3
 2.77298326e-08-4.50893805e-12-3.06512867e+04 5.22593738e+01                   4
C7DIONE                 C   7H  12O   2     G    300.00   3500.00  700.00      1
-7.55853446e-01 8.24536112e-02-4.58824663e-05 1.18274998e-08-1.15807938e-12    2
-3.67546790e+04 2.64722470e+01 3.52180348e+00 5.80098574e-02 6.49700629e-06    3
-3.80577122e-08 1.66580678e-11-3.73535509e+04 7.36075806e+00                   4
NC7H14O                 C   7H  14O   1     G    300.00   3500.00 1490.00      1
 1.37609294e+01 4.99379446e-02-2.21152405e-05 4.72010541e-09-3.98160211e-13    2
-3.97917907e+04-4.67908437e+01-7.39181715e+00 1.06723841e-01-7.92822506e-05    3
 3.02981860e-08-4.68978448e-12-3.34882722e+04 6.36941412e+01                   4
NC7H15-OO               C   7H  15O   2     G    300.00   3500.00 1780.00      1
 2.68006152e+01 3.35780853e-02-1.17982170e-05 1.89992203e-09-1.16218708e-13    2
-2.33388922e+04-1.06550440e+02 1.92333985e+00 8.94820750e-02-5.89083207e-05    3
 1.95441556e-08-2.59434140e-12-1.44825822e+04 2.78126032e+01                   4
NC7-QOOH                C   7H  15O   2     G    300.00   3500.00 1800.00      1
 3.67777396e+01 2.43465609e-02-1.65378967e-05 5.22870320e-09-5.85107826e-13    2
-2.84549754e+04-1.65059582e+02-2.87358719e+00 1.12460620e-01-8.99662796e-05    3
 3.24244006e-08-4.36228802e-12-1.41804978e+04 4.95416697e+01                   4
NC7-OOQOOH              C   7H  15O   4     G    300.00   3500.00 1690.00      1
 2.24694085e+01 4.29307053e-02-1.68910139e-05 3.18431015e-09-2.38592377e-13    2
-4.58962945e+04-7.93472490e+01 2.87430484e+00 8.93096489e-02-5.80557567e-05    3
 1.94228675e-08-2.64074583e-12-3.92731495e+04 2.54699091e+01                   4
C7KETONE                C   7H  14O   1     G    300.00   3500.00 1800.00      1
 1.82994298e+01 4.14393545e-02-1.71834126e-05 3.42714182e-09-2.72037255e-13    2
-4.27848812e+04-6.59785963e+01-2.29236446e-01 8.26141684e-02-5.14957575e-05    3
 1.61354177e-08-2.03707557e-12-3.61145614e+04 3.43024108e+01                   4
NC7-OQOOH               C   7H  14O   3     G    300.00   3500.00 1670.00      1
 2.27584102e+01 4.25741299e-02-1.77950039e-05 3.55398810e-09-2.80791893e-13    2
-5.95329649e+04-8.19251538e+01 2.24997349e+00 9.16961340e-02-6.19165645e-05    3
 2.11673855e-08-2.91752804e-12-5.26831470e+04 2.75334094e+01                   4
NC7H15OOH               C   7H  16O   2     G    300.00   3500.00 1790.00      1
 2.73219576e+01 3.55871014e-02-1.24650786e-05 2.00089299e-09-1.21997718e-13    2
-4.84634175e+04-1.12262051e+02 1.16215161e+00 9.40447685e-02-6.14519505e-05    3
 2.02455380e-08-2.67013250e-12-3.90982069e+04 2.91745384e+01                   4
IC8H16O                 C   8H  16O   1     G    300.00   3500.00 1730.00      1
 2.92525380e+01 3.42835375e-02-1.16024168e-05 1.77292188e-09-1.00402141e-13    2
-4.92824089e+04-1.33818804e+02-8.05235809e+00 1.20537632e-01-8.63892043e-05    3
 3.05924932e-08-4.26508008e-12-3.63749148e+04 6.66033676e+01                   4
IC8H17-OO               C   8H  17O   2     G    300.00   3500.00 1600.00      1
 2.43863205e+01 4.79091902e-02-1.96116195e-05 3.85759248e-09-3.01446152e-13    2
-3.51809034e+04-9.31491912e+01-7.10506864e-01 1.10651259e-01-7.84323086e-05    3
 2.83662129e-08-4.13091810e-12-2.71499187e+04 3.97240934e+01                   4
IC8-QOOH                C   8H  17O   2     G    300.00   3500.00 1560.00      1
 2.59202598e+01 4.65574237e-02-1.91478807e-05 3.78861223e-09-2.97861918e-13    2
-2.91331932e+04-1.00455346e+02-9.92411415e-01 1.15564273e-01-8.55006204e-05    3
 3.21444839e-08-4.84207212e-12-2.07364398e+04 4.13504188e+01                   4
IC8T-QOOH               C   8H  17O   2     G    300.00   3500.00 1560.00      1
 2.59202598e+01 4.65574237e-02-1.91478807e-05 3.78861223e-09-2.97861918e-13    2
-2.91331932e+04-1.00455346e+02-9.92411415e-01 1.15564273e-01-8.55006204e-05    3
 3.21444839e-08-4.84207212e-12-2.07364398e+04 4.13504188e+01                   4
IC8-OOQOOH              C   8H  17O   4     G    300.00   3500.00 1710.00      1
 3.48314344e+01 3.98145837e-02-1.43978156e-05 2.42273023e-09-1.57987515e-13    2
-5.01227423e+04-1.45334583e+02 1.76391251e+00 1.17165512e-01-8.22495073e-05    3
 2.88756315e-08-4.02537074e-12-3.88136498e+04 3.19376018e+01                   4
IC8-OQOOH               C   8H  16O   3     G    300.00   3500.00 1770.00      1
 3.33140848e+01 3.48304637e-02-1.19632298e-05 1.85711996e-09-1.07309755e-13    2
-6.88276642e+04-1.40834056e+02 5.55149631e-01 1.08861956e-01-7.47017824e-05    3
 2.54874599e-08-3.44492839e-12-5.72310012e+04 3.59135519e+01                   4
KHDECA                  C  10H  16O   3     G    300.00   3500.00 1460.00      1
 1.16022413e+01 3.57303676e-02-1.34415895e-05 2.50437497e-09-1.89510332e-13    2
-3.63821555e+04-4.98532931e+01-8.02402160e+00 8.95009509e-02-6.86853394e-05    3
 2.77298316e-08-4.50893783e-12-3.06512867e+04 5.22593734e+01                   4
NC10-OQOOH              C  10H  20O   3     G    300.00   3500.00 1650.00      1
 2.99089218e+01 5.87016504e-02-2.37959602e-05 4.63915061e-09-3.59659380e-13    2
-7.07246440e+04-1.14602314e+02 2.87865558e+00 1.24229568e-01-8.33667947e-05    3
 2.87081747e-08-4.00648121e-12-6.18046561e+04 2.93391851e+01                   4
NC12-OQOOH              C  12H  24O   3     G    300.00   3500.00 1800.00      1
 2.89762386e+01 8.51935374e-02-4.32222255e-05 1.03184958e-08-9.52874267e-13    2
-7.66784398e+04-1.07151219e+02 4.95723497e+00 1.38569101e-01-8.77018619e-05    3
 2.67924352e-08-3.24092140e-12-6.80315985e+04 2.28446393e+01                   4
NC16-OQOOH              C  16H  32O   3     G    300.00   3500.00 1690.00      1
 4.88441403e+01 8.47832934e-02-3.17577342e-05 5.56702310e-09-3.82331041e-13    2
-9.50808943e+04-2.07202689e+02 1.75040576e+00 1.96247754e-01-1.30690687e-04    3
 4.45938291e-08-6.15552719e-12-7.91632120e+04 4.47087840e+01                   4
IC16-OQOOH              C  16H  32O   3     G    300.00   3500.00 1590.00      1
 5.03105850e+01 8.85535133e-02-3.63077758e-05 7.13747459e-09-5.56692445e-13    2
-1.01978072e+05-2.30341226e+02-5.93668615e+00 2.30056082e-01-1.69800765e-04    3
 6.31093780e-08-9.35730619e-12-8.40914402e+04 6.71031167e+01                   4
IC12-OQOOH              C  12H  24O   3     G    300.00   3500.00 1800.00      1
 2.89762386e+01 8.51935374e-02-4.32222255e-05 1.03184958e-08-9.52874267e-13    2
-7.66784398e+04-1.07151219e+02 4.95723497e+00 1.38569101e-01-8.77018619e-05    3
 2.67924352e-08-3.24092140e-12-6.80315985e+04 2.28446393e+01                   4
RMCYC6-OO               C   7H  13O   2     G    300.00   3500.00 1800.00      1
 2.27624353e+01 3.77290578e-02-1.50512016e-05 2.88934761e-09-2.22140217e-13    2
-2.53740840e+04-9.90983455e+01-6.71698854e+00 1.03238889e-01-6.96427272e-05    3
 2.31084312e-08-3.03034627e-12-1.47614915e+04 6.04504459e+01                   4
MCYC6-QOOH              C   7H  13O   2     G    300.00   3500.00 1800.00      1
 2.93659910e+01 2.65374233e-02-8.30521741e-06 1.12153103e-09-5.23348200e-14    2
-2.28599212e+04-1.33867717e+02-7.82169697e+00 1.09176730e-01-7.71713063e-05    3
 2.66274899e-08-3.59482911e-12-9.47235350e+03 6.73998084e+01                   4
MCYC6T-QOOH             C   7H  13O   2     G    300.00   3500.00 1800.00      1
 2.93659910e+01 2.65374233e-02-8.30521741e-06 1.12153103e-09-5.23348200e-14    2
-2.28599212e+04-1.33867717e+02-7.82169697e+00 1.09176730e-01-7.71713063e-05    3
 2.66274899e-08-3.59482911e-12-9.47235350e+03 6.73998084e+01                   4
MCYC6T-OOQOOH           C   7H  13O   4     G    300.00   3500.00 1770.00      1
 3.14587712e+01 3.12961290e-02-1.06604066e-05 1.62769033e-09-9.15069237e-14    2
-4.08526709e+04-1.40718370e+02-4.29317157e+00 1.12091480e-01-7.91310429e-05    3
 2.74170072e-08-3.73406581e-12-2.81964831e+04 5.21777155e+01                   4
MCYC6-OOQOOH            C   7H  13O   4     G    300.00   3500.00 1770.00      1
 3.14587712e+01 3.12961290e-02-1.06604066e-05 1.62769033e-09-9.15069237e-14    2
-4.08526709e+04-1.40718370e+02-4.29317157e+00 1.12091480e-01-7.91310429e-05    3
 2.74170072e-08-3.73406581e-12-2.81964831e+04 5.21777155e+01                   4
KMCYC6                  C   7H  12O   3     G    300.00   3500.00 1800.00      1
 2.89245694e+01 2.89702916e-02-1.00807607e-05 1.60861901e-09-9.81382707e-14    2
-5.92858032e+04-1.29605415e+02-5.14358426e+00 1.04677300e-01-7.31699341e-05    3
 2.49749795e-08-3.34346612e-12-4.70212679e+04 5.47785393e+01                   4
QDECOOH                 C  10H  17O   2     G    300.00   3500.00 1800.00      1
 1.72379170e+01 3.76978752e-02-1.66331319e-05 3.54555193e-09-3.00284997e-13    2
-1.92027470e+04-7.01676441e+01-6.00367530e+00 8.93458581e-02-5.96731176e-05    3
 1.94862874e-08-2.51427603e-12-1.08357738e+04 5.56207018e+01                   4
RDECOO                  C  10H  17O   2     G    300.00   3500.00 1800.00      1
 1.72379170e+01 3.76978752e-02-1.66331319e-05 3.54555193e-09-3.00284997e-13    2
-1.92027470e+04-7.01676441e+01-6.00367530e+00 8.93458581e-02-5.96731176e-05    3
 1.94862874e-08-2.51427603e-12-1.08357738e+04 5.56207018e+01                   4
ZDECA                   C  10H  17O   4     G    300.00   3500.00 1800.00      1
 1.72379170e+01 3.76978752e-02-1.66331319e-05 3.54555193e-09-3.00284997e-13    2
-1.92027470e+04-7.01676441e+01-6.00367530e+00 8.93458581e-02-5.96731176e-05    3
 1.94862874e-08-2.51427603e-12-1.08357738e+04 5.56207018e+01                   4
DECA_ET                 C  10H  16O   1     G    300.00   3500.00 1450.00      1
 2.11071726e+01 5.53253979e-02-2.30739157e-05 4.67748849e-09-3.78388476e-13    2
-3.67326427e+04-9.38585002e+01-2.77500526e+01 1.90103950e-01-1.62500004e-04    3
 6.87814372e-08-1.14307934e-11-2.25640474e+04 1.60002934e+02                   4
NC10H21-OO              C  10H  21O   2     G    300.00   3500.00 1800.00      1
 3.23779961e+01 5.24885097e-02-1.93369945e-05 3.35369138e-09-2.28448249e-13    2
-4.06447326e+04-1.32099033e+02 1.67478092e+00 1.20717877e-01-7.61948004e-05    3
 2.44121380e-08-3.15323250e-12-2.95915751e+04 3.40731730e+01                   4
NC10-QOOH               C  10H  21O   2     G    300.00   3500.00 1800.00      1
 3.67714457e+01 4.56787362e-02-1.56929360e-05 2.49979572e-09-1.53467622e-13    2
-3.72897383e+04-1.54708940e+02 8.46534301e-01 1.25511873e-01-8.22205498e-05    3
 2.71396527e-08-3.57566998e-12-2.43567702e+04 3.97241754e+01                   4
NC10-OOQOOH             C  10H  21O   4     G    300.00   3500.00 1800.00      1
 4.08087612e+01 4.96339769e-02-1.81420284e-05 3.12007174e-09-2.11176095e-13    2
-5.65432917e+04-1.73810959e+02 2.62701411e+00 1.34482304e-01-8.88489674e-05    3
 2.93078269e-08-3.84836432e-12-4.27978628e+04 3.28366210e+01                   4
RODECOO                 C  10H  17O   2     G    300.00   3500.00 1800.00      1
 1.72379170e+01 3.76978752e-02-1.66331319e-05 3.54555193e-09-3.00284997e-13    2
-1.92027470e+04-7.01676441e+01-6.00367530e+00 8.93458581e-02-5.96731176e-05    3
 1.94862874e-08-2.51427603e-12-1.08357738e+04 5.56207018e+01                   4
NC12-QOOH               C  12H  25O   2     G    300.00   3500.00 1800.00      1
 4.28763876e+01 5.51011342e-02-1.90602370e-05 3.05790955e-09-1.89216926e-13    2
-4.53974042e+04-1.84606533e+02 5.27388171e-01 1.49210022e-01-9.74843100e-05    3
 3.21038625e-08-4.22337706e-12-3.01517644e+04 4.45950862e+01                   4
NC12H25-OO              C  12H  25O   2     G    300.00   3500.00 1800.00      1
 3.82754161e+01 6.23046040e-02-2.29785807e-05 3.99220512e-09-2.72630492e-13    2
-4.86703029e+04-1.60846129e+02 1.39669299e+00 1.44257322e-01-9.12725124e-05    3
 2.92862539e-08-3.78569282e-12-3.53939626e+04 3.87492141e+01                   4
NC12-OOQOOH             C  12H  25O   4     G    300.00   3500.00 1800.00      1
 4.68889891e+01 5.84439248e-02-2.09491280e-05 3.49896761e-09-2.27324087e-13    2
-6.45487958e+04-2.03262229e+02 2.75932157e+00 1.56509853e-01-1.02670734e-04    3
 3.37662293e-08-4.43111043e-12-4.86621155e+04 3.55767374e+01                   4
QODECOOH                C  10H  17O   2     G    300.00   3500.00 1800.00      1
 1.72379170e+01 3.76978752e-02-1.66331319e-05 3.54555193e-09-3.00284997e-13    2
-1.92027470e+04-7.01676441e+01-6.00367530e+00 8.93458581e-02-5.96731176e-05    3
 1.94862874e-08-2.51427603e-12-1.08357738e+04 5.56207018e+01                   4
IC12-QOOH               C  12H  25O   2     G    300.00   3500.00 1800.00      1
 4.28763876e+01 5.51011342e-02-1.90602370e-05 3.05790955e-09-1.89216926e-13    2
-4.53974042e+04-1.84606533e+02 5.27388171e-01 1.49210022e-01-9.74843100e-05    3
 3.21038625e-08-4.22337706e-12-3.01517644e+04 4.45950862e+01                   4
IC12H25-OO              C  12H  25O   2     G    300.00   3500.00 1800.00      1
 3.82754161e+01 6.23046040e-02-2.29785807e-05 3.99220512e-09-2.72630492e-13    2
-4.86703029e+04-1.60846129e+02 1.39669299e+00 1.44257322e-01-9.12725124e-05    3
 2.92862539e-08-3.78569282e-12-3.53939626e+04 3.87492141e+01                   4
IC12-OOQOOH             C  12H  25O   4     G    300.00   3500.00 1800.00      1
 4.68889891e+01 5.84439248e-02-2.09491280e-05 3.49896761e-09-2.27324087e-13    2
-6.45487958e+04-2.03262229e+02 2.75932157e+00 1.56509853e-01-1.02670734e-04    3
 3.37662293e-08-4.43111043e-12-4.86621155e+04 3.55767374e+01                   4
NC16H33-OO              C  16H  33O   2     G    300.00   3500.00 1800.00      1
 5.00344411e+01 8.20070293e-02-3.03043085e-05 5.28016955e-09-3.62023094e-13    2
-6.47045844e+04-2.18137165e+02 8.65097451e-01 1.91272237e-01-1.21358649e-04    3
 3.90039992e-08-5.04588833e-12-4.70036207e+04 4.79775805e+01                   4
IC16H33-OO              C  16H  33O   2     G    300.00   3500.00 1460.00      1
 3.94749832e+01 1.06211465e-01-4.74108350e-05 1.02029331e-08-8.67106968e-13    2
-6.81954478e+04-1.73182742e+02-7.55515825e+00 2.35061168e-01-1.79790666e-04    3
 7.06503448e-08-1.12176912e-11-5.44626465e+04 7.15084240e+01                   4
IC16-QOOH               C  16H  33O   2     G    300.00   3500.00 1460.00      1
 4.22439777e+01 1.02589729e-01-4.54459563e-05 9.70909219e-09-8.19910985e-13    2
-6.26654633e+04-1.86283131e+02-7.79323361e+00 2.39677980e-01-1.86290049e-04    3
 7.40214632e-08-1.18323033e-11-4.80545976e+04 7.40533931e+01                   4
IC16T-QOOH              C  16H  33O   2     G    300.00   3500.00 1560.00      1
 5.03537423e+01 8.72534961e-02-3.55849715e-05 6.99644148e-09-5.47406484e-13    2
-6.86133969e+04-2.32227105e+02-7.33743207e+00 2.35179584e-01-1.77821595e-04    3
 6.77813231e-08-1.02885734e-11-5.06137505e+04 7.17539094e+01                   4
NC16-QOOH               C  16H  33O   2     G    300.00   3500.00 1800.00      1
 5.49634958e+01 7.74661646e-02-2.71265545e-05 4.36952893e-09-2.68718580e-13    2
-8.49949322e+04-2.46826109e+02 8.02820430e-02 1.99428862e-01-1.28762136e-04    3
 4.20123367e-08-5.49688633e-12-6.52369753e+04 5.02132937e+01                   4
NC16-OOQOOH             C  16H  33O   4     G    300.00   3500.00 1800.00      1
 5.83925874e+01 7.87490384e-02-2.86987295e-05 4.90944156e-09-3.29403472e-13    2
-8.05061522e+04-2.59208996e+02 2.14519072e+00 2.03743253e-01-1.32860575e-04    3
 4.34879029e-08-5.68752311e-12-6.02570894e+04 4.52136486e+01                   4
IC16-OOQOOH             C  16H  33O   4     G    300.00   3500.00 1420.00      1
 4.21122153e+01 1.11834112e-01-5.11978395e-05 1.12541431e-08-9.72533672e-13    2
-7.89343510e+04-1.80495591e+02-6.54289858e+00 2.48890771e-01-1.95976000e-04    3
 7.92251105e-08-1.29392533e-11-6.51162987e+04 7.12984583e+01                   4
IC16T-OOQOOH            C  16H  33O   4     G    300.00   3500.00 1370.00      1
 4.07769136e+01 1.15135964e-01-5.36319072e-05 1.19826896e-08-1.04989864e-12    2
-8.16821247e+04-1.74509335e+02-7.08781201e+00 2.54886987e-01-2.06643977e-04    3
 8.64411178e-08-1.46372030e-11-6.85671899e+04 7.14786272e+01                   4
RC6H5C4H8OO             C  10H  13O   2     G    300.00   3500.00 1800.00      1
 2.95255354e+01 3.88781195e-02-1.67600168e-05 3.28863964e-09-2.50060931e-13    2
-1.12745934e+04-1.27907214e+02-2.97080496e+00 1.11092209e-01-7.69384248e-05    3
 2.55769389e-08-3.34565805e-12 4.24089083e+02 4.79697592e+01                   4
QC6H5C4H8               C  10H  13O   2     G    300.00   3500.00 1600.00      1
 2.58642212e+01 4.31466573e-02-1.79342318e-05 3.56441946e-09-2.80425987e-13    2
-2.83087866e+03-1.02550355e+02-4.02896128e+00 1.17879613e-01-8.79963783e-05    3
 3.27569805e-08-4.84176364e-12 6.73493973e+03 5.57168746e+01                   4
QC6H5C4H8OO             C  10H  13O   4     G    300.00   3500.00 1340.00      1
 2.21297428e+01 5.89831635e-02-2.79882014e-05 6.34013528e-09-5.60973844e-13    2
-1.94753096e+04-7.75039160e+01-3.35040485e+00 1.35043306e-01-1.13130152e-04    3
 4.86993146e-08-8.46380580e-12-1.26466300e+04 5.28803326e+01                   4
KETBBZ                  C  10H  12O   3     G    300.00   3500.00 1370.00      1
 2.04509776e+01 5.51768872e-02-2.63136967e-05 5.98071120e-09-5.30329154e-13    2
-7.66936916e+03-7.18793093e+01-2.50633155e+00 1.22205527e-01-9.97027184e-05    3
 4.16931305e-08-7.04719399e-12-1.37906645e+03 4.61036442e+01                   4
NC3H7OH                 C   3H   8O   1     G    300.00   3500.00 1800.00      1
 1.10496314e+01 1.81260739e-02-6.48607662e-06 1.10352527e-09-7.45033831e-14    2
-3.64580963e+04-3.27312831e+01-2.51644390e-01 4.32400202e-02-2.74143652e-05    3
 8.85474326e-09-1.15106144e-12-3.23896370e+04 2.84335792e+01                   4
CH3CHCH2OH              C   3H   7O   1     G    300.00   3500.00 1800.00      1
 7.63374910e+00 2.08880280e-02-8.76973957e-06 1.80199698e-09-1.48383965e-13    2
-1.08851845e+04-1.05293328e+01 2.18301323e+00 3.30007744e-02-1.88636949e-05    3
 5.54049896e-09-6.67620350e-13-8.92291954e+03 1.89711868e+01                   4
CH3CH2CHOH              C   3H   7O   1     G    300.00   3500.00 1800.00      1
 1.06992305e+01 1.62004096e-02-6.03307446e-06 1.08995984e-09-7.93898434e-14    2
-1.44167386e+04-2.94436078e+01 9.48802479e-01 3.78680274e-02-2.40894226e-05    3
 7.77749619e-09-1.00821434e-12-1.09065845e+04 2.33277426e+01                   4
CH2CH2CH2OH             C   3H   7O   1     G    300.00   3500.00 1800.00      1
 1.10024647e+01 1.50905463e-02-5.07771848e-06 7.82747443e-10-4.56159339e-14    2
-1.15495010e+04-2.90815210e+01 2.77594430e-01 3.89235913e-02-2.49385893e-05    3
 8.13862553e-09-1.06726567e-12-7.68854770e+03 2.89637141e+01                   4
CH3CH2CH2O              C   3H   7O   1     G    300.00   3500.00 1800.00      1
 6.66433619e+00 2.45624456e-02-1.14187469e-05 2.58003148e-09-2.29895655e-13    2
-7.91390221e+03-8.44864803e+00 1.62185675e+00 3.57679554e-02-2.07566718e-05    3
 6.03852218e-09-7.10241585e-13-6.09860961e+03 1.88423026e+01                   4
IC3H7OH                 C   3H   8O   1     G    300.00   3500.00 1490.00      1
 1.02736704e+01 1.89903304e-02-6.50928475e-06 9.85863113e-10-5.35100946e-14    2
-3.77812750e+04-2.92304764e+01-1.25951107e+00 4.99518914e-02-3.76786414e-05    3
 1.49318840e-08-2.39344649e-12-3.43443869e+04 3.10096147e+01                   4
CH2CHOHCH3              C   3H   7O   1     G    300.00   3500.00 1380.00      1
 6.32694399e+00 2.38762498e-02-1.07376184e-05 2.33737051e-09-2.01069490e-13    2
-1.14217375e+04-3.95690338e+00 6.40756980e-01 4.03579512e-02-2.86525113e-05    3
 1.09919081e-08-1.76892051e-12-9.85234986e+03 2.53070890e+01                   4
CH3COHCH3               C   3H   7O   1     G    300.00   3500.00 1270.00      1
 6.71652559e+00 2.35306503e-02-1.06144751e-05 2.31761640e-09-1.99886335e-13    2
-1.44175085e+04-7.90476225e+00 1.21649825e+00 4.08535711e-02-3.10746177e-05    3
 1.30578488e-08-2.31410530e-12-1.30205016e+04 1.99442898e+01                   4
C3H7CHO                 C   4H   8O   1     G    300.00   3500.00  700.00      1
-9.77279369e-01 5.24983746e-02-3.09762336e-05 8.32680249e-09-8.38156518e-13    2
-2.70767712e+04 3.27194909e+01 3.71554473e+00 2.56822369e-02 2.64869186e-05    3
-4.64000091e-08 1.87071333e-11-2.77337666e+04 1.17531401e+01                   4
RALD4X                  C   4H   7O   1     G    300.00   3500.00 1140.00      1
-3.84911260e+00 5.11968673e-02-2.73583541e-05 6.64027845e-09-6.13455732e-13    2
-5.69209145e+03 4.92440542e+01 6.06312502e+00 1.64170862e-02 1.84045158e-05    3
-2.01216338e-08 5.25538467e-12-7.95208162e+03 1.24454237e-01                   4
C3H5CHO                 C   4H   6O   1     G    300.00   3500.00 1610.00      1
 9.36564374e+00 1.99394665e-02-8.24714101e-06 1.63840860e-09-1.29181838e-13    2
-1.44293666e+04-2.07054062e+01 2.40474632e-01 4.26106940e-02-2.93694027e-05    3
 1.03846868e-08-1.48729956e-12-1.14910622e+04 2.76639773e+01                   4
IC3H5CHO                C   4H   6O   1     G    300.00   3500.00 1370.00      1
 8.96605739e+00 2.20962390e-02-1.00901149e-05 2.22139290e-09-1.91792276e-13    2
-1.79920101e+04-2.11939228e+01 6.92942029e-01 4.62513203e-02-3.65372842e-05    3
 1.50910617e-08-2.54027198e-12-1.57251765e+04 2.13235421e+01                   4
NC4H7OH                 C   4H   8O   1     G    300.00   3500.00 1260.00      1
 9.47752990e+00 2.59932946e-02-1.14395829e-05 2.45196152e-09-2.08596712e-13    2
-2.58308659e+04-2.26233204e+01-1.20059157e+00 5.98920930e-02-5.17952952e-05    3
 2.38041903e-08-4.44515003e-12-2.31399793e+04 3.13602822e+01                   4
IC4H7OH                 C   4H   8O   1     G    300.00   3500.00 1800.00      1
 1.15391972e+01 2.16392208e-02-8.55965895e-06 1.65851695e-09-1.29717210e-13    2
-2.50645504e+04-3.36073962e+01 1.41746548e+00 4.41319580e-02-2.73036066e-05    3
 8.60071980e-09-1.09391205e-12-2.14207270e+04 2.11735275e+01                   4
IC3H7CHO                C   4H   8O   1     G    300.00   3500.00 1800.00      1
 1.25375030e+01 2.06759847e-02-7.90606758e-06 1.44761626e-09-1.05776601e-13    2
-3.22363631e+04-4.10505155e+01-3.44731979e-01 4.93031735e-02-3.17620582e-05    3
 1.02831683e-08-1.33293661e-12-2.75987585e+04 2.86708273e+01                   4
RIBALDB                 C   4H   7O   1     G    300.00   3500.00 1090.00      1
 7.80130141e+00 2.08311675e-02-4.31906608e-06-1.13870025e-10 8.81387193e-14    2
-1.58031223e+03-1.28298252e+01-1.99174488e+00 5.67689520e-02-5.37747329e-05    3
 3.01342442e-08-6.84950216e-12 5.54571864e+02 3.52599044e+01                   4
RIBALDG                 C   4H   7O   1     G    300.00   3500.00 1050.00      1
 9.00440169e+00 1.88029637e-02-3.43463831e-06-2.58096232e-10 9.53220741e-14    2
-4.96767966e+03-1.61872933e+01-3.42297333e+00 6.61453447e-02-7.10666112e-05    3
 4.26828389e-08-1.01287101e-11-2.35793090e+03 4.43739412e+01                   4
N1C4H9OH                C   4H  10O   1     G    300.00   3500.00 1800.00      1
 1.48230800e+01 2.16832750e-02-7.46704059e-06 1.19388933e-09-7.36745605e-14    2
-4.08306214e+04-5.15940710e+01-4.78997507e-01 5.56878917e-02-3.58042211e-05    3
 1.16891414e-08-1.53134846e-12-3.53218735e+04 3.12239646e+01                   4
CH3CH2CHCH2OH           C   4H   9O   1     G    300.00   3500.00 1800.00      1
 1.13530984e+01 2.45578868e-02-9.82948597e-06 1.91527527e-09-1.49940479e-13    2
-1.52382169e+04-2.90980448e+01 1.95582518e+00 4.54407163e-02-2.72318438e-05    3
 8.36059300e-09-1.04512350e-12-1.18551985e+04 2.17619584e+01                   4
CH2CH2CH2CH2OH          C   4H   9O   1     G    300.00   3500.00 1790.00      1
 1.44669861e+01 1.91857582e-02-6.39892818e-06 9.65852380e-10-5.40085895e-14    2
-1.57844516e+04-4.62017114e+01 4.01249151e-02 5.14245541e-02-3.34146789e-05    3
 1.10275845e-08-1.45927844e-12-1.06196353e+04 3.17990982e+01                   4
CH3CH2CH2CH2O           C   4H   9O   1     G    300.00   3500.00 1800.00      1
 9.76394478e+00 2.97115880e-02-1.36105423e-05 3.01462613e-09-2.63554844e-13    2
-1.20864798e+04-2.37714390e+01 1.13482584e+00 4.88874078e-02-2.95903922e-05    3
 8.93308905e-09-1.08556358e-12-8.97999697e+03 2.29311529e+01                   4
CH3CH2CH2CHOH           C   4H   9O   1     G    300.00   3500.00 1800.00      1
 1.45806715e+01 1.95400775e-02-6.85981501e-06 1.13500377e-09-7.38189229e-14    2
-1.88304393e+04-4.88995913e+01 7.07705093e-01 5.03688917e-02-3.25504935e-05    3
 1.06500699e-08-1.39535588e-12-1.38361714e+04 2.61837970e+01                   4
CH3CHCH2CH2OH           C   4H   9O   1     G    300.00   3500.00 1800.00      1
 1.10473988e+01 2.49495901e-02-1.02454978e-05 2.07975683e-09-1.70768002e-13    2
-1.60937894e+04-2.75546714e+01-8.85954576e-02 4.96962441e-02-3.08677094e-05    3
 9.71761299e-09-1.23158136e-12-1.20848314e+04 3.27156527e+01                   4
N2C4H9OH                C   4H  10O   1     G    300.00   3500.00 1800.00      1
 1.39850058e+01 2.35768255e-02-8.73106342e-06 1.51546230e-09-1.02847526e-13    2
-4.24053992e+04-4.83702752e+01 1.11913127e-01 5.44059202e-02-3.44219757e-05    3
 1.10306150e-08-1.42439651e-12-3.74110858e+04 2.67137962e+01                   4
CH2CH2CHOHCH3           C   4H   9O   1     G    300.00   3500.00 1800.00      1
 1.39333099e+01 2.07599762e-02-7.56097133e-06 1.27900106e-09-8.37238451e-14    2
-1.74897437e+04-4.46134923e+01 9.11732959e-01 4.96968138e-02-3.16750027e-05    3
 1.02101238e-08-1.32415756e-12-1.28019760e+04 2.58619985e+01                   4
CH3CH2CHOHCH2           C   4H   9O   1     G    300.00   3500.00 1800.00      1
 1.39333099e+01 2.07599762e-02-7.56097133e-06 1.27900106e-09-8.37238451e-14    2
-1.74897437e+04-4.46134923e+01 9.11732959e-01 4.96968138e-02-3.16750027e-05    3
 1.02101238e-08-1.32415756e-12-1.28019760e+04 2.58619985e+01                   4
CH3CHCHOHCH3            C   4H   9O   1     G    300.00   3500.00 1800.00      1
 1.11523992e+01 2.52912429e-02-1.05179521e-05 2.12392751e-09-1.71553115e-13    2
-1.78095401e+04-2.94209584e+01 6.76902557e-01 4.85701242e-02-2.99170199e-05    3
 9.30876742e-09-1.16944755e-12-1.40383613e+04 2.72746145e+01                   4
CH3CH2COHCH3            C   4H   9O   1     G    300.00   3500.00 1430.00      1
 8.72382313e+00 3.04342821e-02-1.39185542e-05 3.06043840e-09-2.64689208e-13    2
-1.80661274e+04-1.71435120e+01 1.27395826e+00 5.12730649e-02-3.57774173e-05    3
 1.32510506e-08-2.04626476e-12-1.59354661e+04 2.14624058e+01                   4
TC4H9OH                 C   4H  10O   1     G    300.00   3500.00 1440.00      1
 9.08150395e+00 3.22201835e-02-1.41979350e-05 3.03249258e-09-2.56658350e-13    2
-4.23917231e+04-2.36263222e+01-6.99999550e-01 5.93910265e-02-4.25008965e-05    3
 1.61357155e-08-2.53152344e-12-3.95746501e+04 2.71305358e+01                   4
RTC4H8OH                C   4H   9O   1     G    300.00   3500.00 1380.00      1
 8.66823606e+00 3.01271702e-02-1.35256231e-05 2.94117221e-09-2.52822111e-13    2
-1.73478970e+04-1.68023785e+01 1.39880725e-03 5.52484376e-02-4.08313485e-05    3
 1.61323439e-08-2.64252713e-12-1.49558499e+04 2.78015466e+01                   4
IC4H9OH                 C   4H  10O   1     G    300.00   3500.00 1800.00      1
 1.44537508e+01 2.20810711e-02-7.57959413e-06 1.19533698e-09-7.16167878e-14    2
-4.15822807e+04-5.13315448e+01-5.45479347e-01 5.54126937e-02-3.53559463e-05    3
 1.14828748e-08-1.50044149e-12-3.61825578e+04 2.98474178e+01                   4
CH3CHCH3CHOH            C   4H   9O   1     G    300.00   3500.00 1450.00      1
 8.91411937e+00 2.94184828e-02-1.30488491e-05 2.81020917e-09-2.39749766e-13    2
-1.71145337e+04-1.85255728e+01 6.16106295e-01 5.23095533e-02-3.67292669e-05    3
 1.36977576e-08-2.11691329e-12-1.47081099e+04 2.45907828e+01                   4
CH3CCH2OHCH3            C   4H   9O   1     G    300.00   3500.00  700.00      1
 2.02076663e+00 4.09903682e-02-2.06486865e-05 5.00507643e-09-4.71523446e-13    2
-1.40718373e+04 2.15880986e+01 3.53447953e+00 3.23405802e-02-2.11342645e-06    3
-1.26475522e-08 5.83298677e-12-1.42837571e+04 1.48252123e+01                   4
CH2CHCH2OHCH3           C   4H   9O   1     G    300.00   3500.00 1780.00      1
 1.38129862e+01 2.02819149e-02-7.03373606e-06 1.12440102e-09-6.86005419e-14    2
-1.64045558e+04-4.42516768e+01 2.32452984e-01 5.07999670e-02-3.27511957e-05    3
 1.07564084e-08-1.42141056e-12-1.15698860e+04 2.90972624e+01                   4
MEK                     C   4H   8O   1     G    300.00   3500.00 1800.00      1
 1.00996647e+01 2.22850980e-02-8.24113164e-06 1.42760471e-09-9.77655945e-14    2
-3.40270934e+04-2.55002661e+01 1.67138648e+00 4.10146052e-02-2.38490543e-05    3
 7.20831681e-09-9.00642276e-13-3.09929132e+04 2.01153340e+01                   4
C5H9OH                  C   5H  10O   1     G    300.00   3500.00 1210.00      1
 1.31847861e+01 3.05720282e-02-1.32292714e-05 2.77400172e-09-2.30719066e-13    2
-2.99739273e+04-4.19054271e+01-3.87325767e+00 8.69622556e-02-8.31345119e-05    3
 4.12892857e-08-8.18842238e-12-2.58458807e+04 4.36413840e+01                   4
C4H9CHO                 C   5H  10O   1     G    300.00   3500.00  760.00      1
-1.78433167e+00 6.31204384e-02-3.60836197e-05 9.48321915e-09-9.39522539e-13    2
-2.97113509e+04 3.92478706e+01 5.53298991e+00 2.46082195e-02 3.99273386e-05    3
-5.71930600e-08 2.09934640e-11-3.08235838e+04 5.95416644e+00                   4
IC5H9OH                 C   5H  10O   1     G    300.00   3500.00 1340.00      1
 1.04339671e+01 3.43709898e-02-1.53823536e-05 3.33540404e-09-2.86051952e-13    2
-3.01866096e+04-2.68956282e+01-1.89607132e+00 7.11770745e-02-5.65831947e-05    3
 2.38333350e-08-4.11029280e-12-2.68821593e+04 3.61983073e+01                   4
IC4H9CHO                C   5H  10O   1     G    300.00   3500.00 1800.00      1
 1.47934382e+01 2.65660093e-02-1.04284272e-05 1.98344167e-09-1.51387814e-13    2
-3.60342984e+04-5.12505605e+01 7.73443223e-01 5.77215537e-02-3.63913809e-05    3
 1.15993505e-08-1.48693070e-12-3.09871002e+04 2.46285772e+01                   4
RALD5X                  C   5H   9O   1     G    300.00   3500.00  750.00      1
-3.04813036e-01 5.67977502e-02-3.24057644e-05 8.50471990e-09-8.41763295e-13    2
-5.21420511e+03 3.41933258e+01 6.22525319e+00 2.19707304e-02 3.72482754e-05    3
-5.34099821e-08 1.97964707e-11-6.19371505e+03 4.56811396e+00                   4
ALDC6                   C   6H  12O   1     G    300.00   3500.00 1800.00      1
 1.43376052e+01 3.78182963e-02-1.64821906e-05 3.50930001e-09-2.98005839e-13    2
-3.75955825e+04-4.53859613e+01 1.31726263e+00 6.67523909e-02-4.05939361e-05    3
 1.24395761e-08-1.53832196e-12-3.29082592e+04 2.50828488e+01                   4
RALD6X                  C   6H  11O   1     G    300.00   3500.00 1160.00      1
 5.47459318e-01 6.16901251e-02-2.98352979e-05 6.64392100e-09-5.73135835e-13    2
-1.27523068e+04 2.98980233e+01 4.05975344e+00 4.95787661e-02-1.41740577e-05    3
-2.35679173e-09 1.36667294e-12-1.35671590e+04 1.24319397e+01                   4
C5H11OH                 C   5H  12O   1     G    300.00   3500.00 1800.00      1
 1.84921326e+01 2.54356027e-02-8.57802765e-06 1.32118770e-09-7.66434680e-14    2
-4.51605170e+04-6.98750070e+01-6.77484565e-01 6.80347520e-02-4.40773187e-05    3
 1.44690733e-08-1.90273869e-12-3.82594548e+04 3.38749602e+01                   4
RPENT1OHA               C   5H  11O   1     G    300.00   3500.00 1800.00      1
 1.84065772e+01 2.29900187e-02-7.76357340e-06 1.20244130e-09-7.05741205e-14    2
-2.32226149e+04-6.80495345e+01 4.75636978e-01 6.28365525e-02-4.09690182e-05    3
 1.35007542e-08-1.77867313e-12-1.67674764e+04 2.89964545e+01                   4
RPENT1OHB               C   5H  11O   1     G    300.00   3500.00 1800.00      1
 1.50707238e+01 2.82315413e-02-1.08918043e-05 2.02927062e-09-1.51568824e-13    2
-1.95906720e+04-4.76575400e+01 1.72826110e+00 5.78814583e-02-3.56000685e-05    3
 1.11804796e-08-1.42257007e-12-1.47873854e+04 2.45546514e+01                   4
IC5H11OH                C   5H  12O   1     G    300.00   3500.00 1800.00      1
 1.75261752e+01 2.67328609e-02-9.21963365e-06 1.46159055e-09-8.81570173e-14    2
-4.58408775e+04-6.62686630e+01-6.91391533e-01 6.72163424e-02-4.29558683e-05    3
 1.39564923e-08-1.82356003e-12-3.92825534e+04 3.23286084e+01                   4
RIPENTOHA               C   5H  11O   1     G    300.00   3500.00 1620.00      1
 1.36179093e+01 3.09491084e-02-1.25439327e-05 2.45214985e-09-1.90908922e-13    2
-2.20274845e+04-4.25086925e+01 6.58084951e-01 6.29486746e-02-4.21731607e-05    3
 1.46452478e-08-2.07255984e-12-1.78285014e+04 2.62671266e+01                   4
RIPENTOHB               C   5H  11O   1     G    300.00   3500.00 1800.00      1
 1.43827461e+01 2.99341331e-02-1.24371790e-05 2.55512971e-09-2.11814040e-13    2
-2.12442488e+04-4.60019589e+01-6.44589008e-01 6.33282112e-02-4.02655775e-05    3
 1.28619439e-08-1.64331602e-12-1.58344082e+04 3.53291137e+01                   4
C6H13OH                 C   6H  14O   1     G    300.00   3500.00 1800.00      1
 2.78613505e+01 1.77437757e-02-2.99502444e-06 1.18963293e-11 2.84574013e-14    2
-5.19282562e+04-1.19896997e+02-1.83303812e+00 8.37313060e-02-5.79846331e-05    3
 2.03784180e-08-2.80022617e-12-4.12382763e+04 4.08152287e+01                   4
RHEX1OHA                C   6H  13O   1     G    300.00   3500.00 1800.00      1
 2.84298221e+01 1.33218221e-02-9.68172392e-07-3.32584677e-10 4.90834902e-14    2
-3.02913851e+04-1.20327872e+02-1.87679993e-01 7.69162711e-02-5.39635466e-05    3
 1.92953317e-08-2.67701600e-12-1.99890844e+04 3.45560186e+01                   4
RHEX1OHB                C   6H  13O   1     G    300.00   3500.00 1800.00      1
 2.97416429e+01 1.08284393e-02 6.26458164e-07-7.76125681e-10 9.43842379e-14    2
-2.87904782e+04-1.27477420e+02-8.09485813e-02 7.71008648e-02-5.46005631e-05    3
 1.96783266e-08-2.74651192e-12-1.80543453e+04 3.39286666e+01                   4
NC5H12                  C   5H  12          G    300.00   3500.00 1800.00      1
 2.12559079e+01 1.49866380e-02-1.56738349e-06-4.84518332e-10 9.00436406e-14    2
-2.80668701e+04-9.05497656e+01-1.97000861e+00 6.65997859e-02-4.45783401e-05    3
 1.54454656e-08-2.12245413e-12-1.97055401e+04 3.51537399e+01                   4
NC5H11                  C   5H  11          G    300.00   3500.00 1800.00      1
 6.93194096e+00 3.75440926e-02-1.65478525e-05 3.53633529e-09-2.99976587e-13    2
-1.73087194e+03-8.88712387e+00-3.57520480e+00 6.08933054e-02-3.60055299e-05    3
 1.07428825e-08-1.30088592e-12 2.05170053e+03 4.79797409e+01                   4
NEOC5H12                C   5H  12          G    300.00   3500.00 1700.00      1
 1.58220754e+01 2.73824194e-02-1.01392663e-05 1.77707245e-09-1.22757215e-13    2
-2.85196990e+04-6.62488213e+01-2.62463400e+00 7.07864416e-02-4.84369329e-05    3
 1.67957652e-08-2.33138851e-12-2.22478178e+04 3.25342335e+01                   4
NEOC5H11                C   5H  11          G    300.00   3500.00 1670.00      1
 1.43276271e+01 2.66845614e-02-1.02158290e-05 1.86929181e-09-1.35803393e-13    2
-2.94216357e+03-5.15145674e+01-1.29689692e+00 6.41085711e-02-4.38302090e-05    3
 1.52882060e-08-2.14462288e-12 2.27642746e+03 3.18773544e+01                   4
NC5H10                  C   5H  10          G    300.00   3500.00 1800.00      1
 1.11929688e+01 2.82582319e-02-1.13863907e-05 2.22526679e-09-1.74281184e-13    2
-1.02483424e+04-3.39253269e+01-6.89551558e-01 5.46638328e-02-3.33910581e-05    3
 1.03751436e-08-1.30620852e-12-5.97063508e+03 3.03853523e+01                   4
NC5H9-3                 C   5H   9          G    300.00   3500.00 1800.00      1
 9.88286994e+00 2.86275431e-02-1.23662483e-05 2.58308667e-09-2.14521125e-13    2
 7.14211786e+03-2.81379541e+01-9.61360365e-01 5.27258326e-02-3.24481563e-05    3
 1.00208304e-08-1.24754108e-12 1.10460408e+04 3.05532826e+01                   4
B1M2                    C   5H  10          G    300.00   3500.00 1800.00      1
 1.21299360e+01 2.65376107e-02-1.02995501e-05 1.93064471e-09-1.45051143e-13    2
-1.11266099e+04-3.96207308e+01-6.39002261e-01 5.49130291e-02-3.39457321e-05    3
 1.06884899e-08-1.36141853e-12-6.52979208e+03 2.94874270e+01                   4
B1M3                    C   5H  10          G    300.00   3500.00 1800.00      1
 1.31681355e+01 2.49963308e-02-9.30063248e-06 1.64277897e-09-1.14892394e-13    2
-1.09953806e+04-4.60629075e+01-8.44094847e-01 5.61346205e-02-3.52492072e-05    3
 1.12533622e-08-1.44969562e-12-5.95097767e+03 2.97742064e+01                   4
B2M2                    C   5H  10          G    300.00   3500.00 1800.00      1
 9.73411455e+00 3.08235277e-02-1.30973032e-05 2.71635525e-09-2.25270538e-13    2
-1.14704805e+04-2.74876891e+01 1.14407574e-01 5.22006543e-02-3.09115754e-05    3
 9.31423383e-09-1.14164256e-12-8.00738600e+03 2.45761718e+01                   4
CYC5H8                  C   5H   8          G    300.00   3500.00 1460.00      1
 8.43099926e+00 2.71082711e-02-1.07932860e-05 1.95387658e-09-1.31111165e-13    2
-1.09862541e+03-2.37608453e+01-6.56863981e+00 6.82031727e-02-5.30140752e-05    3
 2.12327758e-08-3.43229254e-12 3.28126920e+03 5.42801525e+01                   4
C5H7                    C   5H   7          G    300.00   3500.00 1430.00      1
 7.72404439e+00 2.56072217e-02-8.76350476e-06 8.66194459e-10 3.30416101e-14    2
 2.30808144e+04-1.69352889e+01 2.31765187e-01 4.65646460e-02-3.07468170e-05    3
 1.11148249e-08-1.75867700e-12 2.52236063e+04 2.18904241e+01                   4
LC5H8                   C   5H   8          G    300.00   3500.00 1430.00      1
 8.95829174e+00 2.51033000e-02-8.43679224e-06 8.19905600e-10 3.11426525e-14    2
 4.67953295e+03-2.40439636e+01 1.19183495e+00 4.68276546e-02-3.12245768e-05    3
 1.14435814e-08-1.82614333e-12 6.90073959e+03 1.62025641e+01                   4
DIALLYL                 C   6H  10          G    300.00   3500.00 1670.00      1
 1.46885453e+01 2.58341352e-02-9.34005599e-06 1.60362155e-09-1.08722165e-13    2
 2.72208400e+03-5.11904177e+01-8.93390831e-01 6.31561378e-02-4.28628128e-05    3
 1.49859596e-08-2.11206618e-12 7.92645066e+03 3.19742017e+01                   4
RC6H9A                  C   6H   9          G    300.00   3500.00 1310.00      1
 1.02179197e+01 3.31131701e-02-1.50182304e-05 3.28859670e-09-2.83959245e-13    2
 2.30740211e+04-2.53806634e+01-2.61882183e+00 7.23093274e-02-5.98993265e-05    3
 2.61288492e-08-4.64278605e-12 2.64372474e+04 4.00154625e+01                   4
CYC6H8                  C   6H   8          G    300.00   3500.00 1490.00      1
 8.66772199e+00 3.45074871e-02-1.63846792e-05 3.69261012e-09-3.24421067e-13    2
 5.74022162e+03-2.73566174e+01-6.91358131e+00 7.63364892e-02-5.84944129e-05    3
 2.25336543e-08-3.48567009e-12 1.03834500e+04 5.40276158e+01                   4
CYC6H10                 C   6H  10          G    300.00   3500.00 1800.00      1
 1.51624818e+01 2.76360098e-02-1.05259913e-05 1.89586516e-09-1.35054930e-13    2
-9.29985089e+03-6.25064336e+01-6.01517617e+00 7.46974719e-02-4.97438764e-05    3
 1.64210078e-08-2.15243585e-12-1.67589403e+03 5.21114690e+01                   4
RCYC6H9                 C   6H   9          G    300.00   3500.00 1800.00      1
 1.41670491e+01 2.75651285e-02-1.13337580e-05 2.23021556e-09-1.74683350e-13    2
 7.93866227e+03-5.85442131e+01-6.48639387e+00 7.34616684e-02-4.95808746e-05    3
 1.63958143e-08-2.14212762e-12 1.53739017e+04 5.32365287e+01                   4
CYC6H12                 C   6H  12          G    300.00   3500.00 1800.00      1
 1.12578117e+01 4.34354058e-02-2.02455747e-05 4.54245216e-09-4.01195093e-13    2
-2.30439971e+04-4.47863484e+01-9.43363143e+00 8.94163905e-02-5.85630620e-05    3
 1.87341141e-08-2.37225925e-12-1.55950776e+04 6.72000582e+01                   4
CYC6H11                 C   6H  11          G    300.00   3500.00 1800.00      1
 1.12879146e+01 3.94798452e-02-1.80474797e-05 3.97977166e-09-3.47933742e-13    2
 4.69936135e+02-4.15743397e+01-9.20200331e+00 8.50129960e-02-5.59917721e-05    3
 1.80332133e-08-2.29980063e-12 7.84630657e+03 6.93213702e+01                   4
NC6H12                  C   6H  12          G    300.00   3500.00 1780.00      1
 2.80951656e+01 5.24635940e-03 6.43208126e-06-3.19131383e-09 4.01093690e-13    2
-1.79767848e+04-1.24497293e+02-1.85358323e+00 7.25469185e-02-5.02818730e-05    3
 1.80498675e-08-2.58221830e-12-7.31503023e+03 3.72569570e+01                   4
NC7H16                  C   7H  16          G    300.00   3500.00 1800.00      1
 3.10696108e+01 1.73458885e-02-4.57665256e-07-1.06280927e-09 1.59098821e-13    2
-3.76541587e+04-1.40920491e+02-2.76912798e+00 9.25430859e-02-6.31219964e-05    3
 2.21462023e-08-3.06437500e-12-2.54722127e+04 4.22218224e+01                   4
NC7H15                  C   7H  15          G    300.00   3500.00 1800.00      1
 1.58938328e+01 4.32851136e-02-1.83429559e-05 3.81524521e-09-3.18291849e-13    2
-8.33589320e+03-5.34388041e+01-1.03213633e+00 8.08983783e-02-4.96873431e-05    3
 1.54242775e-08-1.93065745e-12-2.24254432e+03 3.81680717e+01                   4
NC7H14                  C   7H  14          G    300.00   3500.00 1800.00      1
 1.82668066e+01 3.59607967e-02-1.37346455e-05 2.52229198e-09-1.85248391e-13    2
-1.87497330e+04-6.92309052e+01-1.22797275e+00 7.92825285e-02-4.98360887e-05    3
 1.58931969e-08-2.04231851e-12-1.17316124e+04 3.62789074e+01                   4
NC7H13                  C   7H  13          G    300.00   3500.00 1800.00      1
 9.88286994e+00 2.86275431e-02-1.23662483e-05 2.58308667e-09-2.14521125e-13    2
 7.14211786e+03-2.81379541e+01-9.61360365e-01 5.27258326e-02-3.24481563e-05    3
 1.00208304e-08-1.24754108e-12 1.10460408e+04 3.05532826e+01                   4
IC8H18                  C   8H  18          G    300.00   3500.00 1390.00      1
 2.06155889e+01 4.43694084e-02-1.35968850e-05 1.75327596e-09-6.83090585e-14    2
-3.76580615e+04-8.42148814e+01-5.96912086e+00 1.20872170e-01-9.61538223e-05    3
 4.13489294e-08-7.18982946e-12-3.02675122e+04 5.27954204e+01                   4
IC8H17                  C   8H  17          G    300.00   3500.00 1530.00      1
 2.65104236e+01 3.01796800e-02-5.82184855e-06 1.42081429e-11 7.60111260e-14    2
-1.80373027e+04-1.14981200e+02-3.32961206e+00 1.08192845e-01-8.23053437e-05    3
 3.33403498e-08-5.36943686e-12-8.90625183e+03 4.16697269e+01                   4
IC8H16                  C   8H  16          G    300.00   3500.00 1400.00      1
 1.88616064e+01 4.14292809e-02-1.28170534e-05 1.66806697e-09-6.58961250e-14    2
-2.24684067e+04-7.38514304e+01-5.35586566e+00 1.10622058e-01-8.69521720e-05    3
 3.69705044e-08-6.36990281e-12-1.56875145e+04 5.11323804e+01                   4
DIMEPTD                 C   7H  12          G    300.00   3500.00 1310.00      1
 1.53755540e+01 3.27318297e-02-1.05955719e-05 1.52102666e-09-7.69416312e-14    2
-6.19682914e+03-5.37226018e+01-1.29247803e+00 8.36265841e-02-6.88720082e-05    3
 3.11782461e-08-5.73671634e-12-1.82980474e+03 3.11918389e+01                   4
C7H8                    C   7H   8          G    200.00   3500.00 1740.00      1
 1.92535098e+01 1.64137622e-02-3.61136080e-06 2.27428602e-11 5.04456421e-14    2
-3.67626193e+03-8.27561014e+01-4.42382857e+00 7.08444251e-02-5.05343461e-05    3
 1.80008982e-08-2.53262265e-12 4.56345183e+03 4.45878948e+01                   4
C6H5OH                  C   6H   6O   1     G    300.00   3500.00 1330.00      1
 1.39867715e+01 2.02277638e-02-7.36599472e-06 1.21196281e-09-7.46104950e-14    2
-1.80542264e+04-5.08485823e+01-5.47325444e+00 7.87541576e-02-7.33732057e-05    3
 3.42982841e-08-6.29384382e-12-1.28778595e+04 4.85843834e+01                   4
C6H5CHO                 C   7H   6O   1     G    200.00   3500.00 1630.00      1
 2.06104934e+01 1.34209231e-02-2.83635976e-06-5.48104087e-11 5.23167160e-14    2
-1.43315559e+04-8.70895589e+01-3.50845138e+00 7.26085177e-02-5.73034713e-05    3
 2.22221268e-08-3.36439145e-12-6.46877992e+03 4.10544420e+01                   4
C6H5CO                  C   7H   5O   1     G    300.00   3500.00 1470.00      1
 1.31799073e+01 2.42895741e-02-1.09067414e-05 2.35371933e-09-2.00195261e-13    2
 5.86598832e+03-4.37756574e+01-1.56203244e+00 6.44036959e-02-5.18395188e-05    3
 2.09173372e-08-3.35727313e-12 1.02001186e+04 3.30251954e+01                   4
C7H7                    C   7H   7          G    200.00   3500.00 1600.00      1
 1.77148777e+01 1.72901847e-02-4.74309376e-06 3.88421922e-10 1.27959162e-14    2
 1.68881059e+04-7.24712943e+01-3.23806377e+00 6.96725384e-02-5.38515504e-05    3
 2.08502788e-08-3.18436923e-12 2.35930472e+04 3.84624949e+01                   4
CH3C6H4                 C   7H   7          G    200.00   3500.00 1730.00      1
 1.83842194e+01 1.52647323e-02-3.43004161e-06 5.73656533e-11 4.21798590e-14    2
 2.84624019e+04-7.44700991e+01-2.82564606e+00 6.43048837e-02-4.59504041e-05    3
 1.64428618e-08-2.32566640e-12 3.58010154e+04 3.94808227e+01                   4
C6H5O                   H   5C   6O   1     G    100.00   3500.00 1800.00      1
 1.20320201e+01 2.29423294e-02-1.10171048e-05 2.53057349e-09-2.25735875e-13    2
 2.17285930e+02-4.10084397e+01 4.06305261e-01 4.87772513e-02-3.25462064e-05    3
 1.05043148e-08-1.33319994e-12 4.40254327e+03 2.19123542e+01                   4
BENZYNE                 C   6H   4          G    300.00   3500.00 1400.00      1
 1.09465826e+01 1.50373225e-02-5.27844785e-06 8.14607006e-10-4.49072710e-14    2
 5.03301416e+04-3.53782974e+01-3.73796174e+00 5.69931636e-02-5.02311347e-05    3
 2.22206484e-08-3.86741466e-12 5.44418140e+04 4.04070822e+01                   4
RCATEC                  C   6H   5O   2     G    300.00   3500.00 1140.00      1
 1.40810372e+01 2.16036547e-02-9.34848622e-06 1.81734354e-09-1.31737694e-13    2
-2.57458618e+04-4.55416694e+01-4.82568620e+00 8.79430352e-02-9.66371448e-05    3
 5.28633427e-08-1.13260358e-11-2.14351289e+04 4.81496572e+01                   4
C6H4O2                  C   6H   4O   2     G    300.00   3500.00 1410.00      1
 1.74929565e+01 1.29021316e-02-2.02976884e-06-3.72417076e-10 8.59744872e-14    2
-2.22100454e+04-6.49015772e+01-5.23446560e+00 7.73770880e-02-7.06201479e-05    3
 3.20580222e-08-5.66410340e-12-1.58009124e+04 5.25540050e+01                   4
CYC5H4O                 C   5H   4O   1     G    300.00   3500.00 1260.00      1
 6.34459567e+00 2.39841579e-02-8.32755426e-06 8.47127788e-10 2.86249324e-14    2
 3.08659311e+03-9.73181495e+00-5.14379341e+00 6.04552344e-02-5.17455024e-05    3
 2.38195871e-08-4.52940271e-12 5.98166716e+03 4.83481228e+01                   4
C7H7O2                  C   7H   7O   2     G    300.00   3500.00 1420.00      1
 1.76964630e+01 2.58808944e-02-1.00755981e-05 1.78285096e-09-1.17592436e-13    2
 6.43630889e+03-6.45881502e+01-4.45172577e+00 8.82701586e-02-7.59797504e-05    3
 3.27237675e-08-5.56493690e-12 1.27263945e+04 5.00304725e+01                   4
O2C6H4CH3               C   7H   7O   2     G    300.00   3500.00 1300.00      1
 1.57011685e+01 2.91723919e-02-1.27991944e-05 2.73382211e-09-2.31734838e-13    2
 5.63564286e+03-5.46747886e+01-5.21645080e+00 9.35342975e-02-8.70629317e-05    3
 4.08177900e-08-7.55557481e-12 1.10742239e+04 5.17286690e+01                   4
OC6H4CH2                C   7H   6O   1     G    300.00   3500.00 1390.00      1
 1.45795351e+01 2.32519422e-02-8.58329263e-06 1.38947425e-09-7.81466604e-14    2
-5.01093385e+02-5.31869685e+01-4.82277800e+00 7.90859366e-02-6.88358046e-05    3
 3.02875615e-08-5.27564437e-12 4.89274964e+03 4.68072308e+01                   4
C6H5CH2O                C   7H   7O   1     G    300.00   3500.00 1650.00      1
 1.54569212e+01 2.51288554e-02-9.88344503e-06 1.85206287e-09-1.37473897e-13    2
 6.00712904e+03-5.64456921e+01-4.49397746e+00 7.34946703e-02-5.38523676e-05    3
 1.96172841e-08-2.82917408e-12 1.25909256e+04 4.97967780e+01                   4
BZCOOH                  C   7H   8O   2     G    300.00   3500.00 1550.00      1
 1.78036110e+01 3.06807103e-02-1.34555328e-05 2.81495337e-09-2.31878474e-13    2
-1.15055066e+04-6.47324102e+01-3.42659307e+00 8.54683337e-02-6.64758135e-05    3
 2.56193752e-08-3.91001102e-12-4.92414334e+03 4.69952938e+01                   4
C6H5O2                  C   6H   5O   2     G    300.00   3500.00 1300.00      1
 1.17436578e+01 2.50264956e-02-1.11158411e-05 2.39771138e-09-2.04780262e-13    2
 1.03023082e+04-3.29345636e+01-2.98072576e+00 7.03322911e-02-6.33917590e-05    3
 2.92058744e-08-5.36019623e-12 1.41306479e+04 4.19652276e+01                   4
RBBENZ                  C  14H  13          G    300.00   3500.00 1750.00      1
 5.34298817e+01-2.73975002e-03 1.40930443e-05-5.29858171e-09 5.98002314e-13    2
 9.33192483e+03-2.64139632e+02-8.67312012e+00 1.39209969e-01-1.07578143e-04    3
 4.10523468e-08-6.02355890e-12 3.10679755e+04 7.02252737e+01                   4
STILB                   C  14H  12          G    300.00   3500.00 1470.00      1
 3.31295388e+01 3.16424074e-02-7.88066301e-06 4.81368480e-10 4.43951941e-14    2
 1.37146842e+04-1.52659614e+02-1.11031625e+01 1.52003499e-01-1.30698104e-04    3
 5.61808881e-08-9.42831222e-12 2.67190984e+04 7.77787975e+01                   4
OOC6H4OH                H   5C   6O   3     G    100.00   3500.00 1570.00      1
 2.76569235e+01 2.91344224e-04 5.46428566e-06-2.09157809e-09 2.40972818e-13    2
-1.39658762e+04-1.18517528e+02-4.81896333e-01 7.19826049e-02-6.30305493e-05    3
 2.69932775e-08-4.39037362e-12-5.13028675e+03 2.99287474e+01                   4
C6H4OH                  C   6H   5O   1     G    300.00   3500.00 1170.00      1
 1.35501568e+01 1.98692214e-02-8.43356568e-06 1.70584566e-09-1.35582605e-13    2
 1.32571077e+04-4.75538985e+01-6.19433362e+00 8.73717527e-02-9.49752725e-05    3
 5.10173595e-08-1.06722309e-11 1.78773184e+04 5.08018133e+01                   4
C7H6                    C   7H   6          G    300.00   3500.00 1290.00      1
 1.11282370e+01 2.73165788e-02-1.25329630e-05 2.76951365e-09-2.40721321e-13    2
 3.69620903e+04-3.50553552e+01-3.97785310e+00 7.41571682e-02-6.69987646e-05    3
 3.09172147e-08-5.69570215e-12 4.08594615e+04 4.16694455e+01                   4
C7H5                    C   7H   5          G    300.00   3500.00 1250.00      1
 1.21079562e+01 2.22665283e-02-9.87308020e-06 2.11666725e-09-1.79360787e-13    2
 5.15977924e+04-3.78517172e+01-2.81419578e+00 7.00174146e-02-6.71741438e-05    3
 3.26772345e-08-6.29147423e-12 5.53283304e+04 3.74688222e+01                   4
CYC5H4                  C   5H   4          G    200.00   3500.00 1310.00      1
 6.52292988e+00 1.75112089e-02-7.24525129e-06 1.36813986e-09-9.77801453e-14    2
 6.01459585e+04-1.09295502e+01-1.67820648e+00 4.25528466e-02-3.59188823e-05    3
 1.59603185e-08-2.88254706e-12 6.22946562e+04 3.08507214e+01                   4
C5H3                    C   5H   3          G    300.00   3500.00 1370.00      1
 1.06729919e+01 9.74586530e-03-3.33881905e-06 5.09387794e-10-2.86889962e-14    2
 6.39774217e+04-2.94129055e+01 3.35962368e+00 3.10987653e-02-2.67179067e-05    3
 1.18860728e-08-2.10472640e-12 6.59812846e+04 8.17219565e+00                   4
C5H2                    C   5H   2          G    300.00   3500.00 1260.00      1
 1.08586493e+01 8.25356602e-03-3.15379484e-06 5.51063259e-10-3.71272549e-14    2
 7.89908994e+04-3.35264716e+01 1.78531798e+00 3.70577925e-02-3.74445407e-05    3
 1.86943150e-08-3.63697880e-12 8.12773789e+04 1.23440605e+01                   4
C5H5O                   C   5H   5O   1     G    300.00   3500.00 1450.00      1
 1.05801391e+01 2.13128782e-02-9.63052925e-06 2.09384795e-09-1.79321200e-13    2
 1.62543411e+04-3.26154739e+01-4.01979399e+00 6.15885557e-02-5.12950232e-05    3
 2.12499371e-08-3.48209519e-12 2.04883217e+04 4.32455667e+01                   4
LC6H6                   C   6H   6          G    300.00   3500.00 1250.00      1
 1.28863873e+01 1.90072469e-02-7.30992638e-06 1.31482522e-09-9.21386108e-14    2
 3.55364843e+04-4.09021919e+01-1.05889388e+00 6.36321467e-02-6.08598062e-05    3
 2.98747611e-08-5.80412579e-12 3.90228046e+04 2.94875283e+01                   4
C6H4C2H3                C   8H   7          G    200.00   3500.00 1580.00      1
 1.99256074e+01 1.67315531e-02-4.18312959e-06 2.15370082e-10 3.07179836e-14    2
 3.89930313e+04-8.19571073e+01-3.96125907e+00 7.72046328e-02-6.15942812e-05    3
 2.44394847e-08-3.80221154e-12 4.65412811e+04 4.42096618e+01                   4
CRESOL                  C   7H   8O   1     G    300.00   3500.00 1310.00      1
 1.22673689e+01 3.34155277e-02-1.38949865e-05 2.56768147e-09-1.71519537e-13    2
-2.17187244e+04-3.95715135e+01-4.41843935e+00 8.43645604e-02-7.22335736e-05    3
 3.22565298e-08-5.83733030e-12-1.73470426e+04 4.54334869e+01                   4
RCRESOLC                C   7H   7O   1     G    300.00   3500.00 1150.00      1
 1.31541707e+01 2.50657194e-02-5.32353956e-06-2.12687447e-10 1.25840443e-13    2
-3.38086414e+03-4.22339543e+01-6.42956802e+00 9.31830715e-02-9.41722596e-05    3
 5.12938170e-08-1.10712257e-11 1.12339577e+03 5.49833259e+01                   4
RCRESOLO                C   7H   7O   1     G    300.00   3500.00 1150.00      1
 1.27824815e+01 2.40796404e-02-4.51347913e-06-4.25076450e-10 1.44988503e-13    2
-3.97704757e+03-4.00543789e+01-6.60757190e+00 9.15233043e-02-9.24834755e-05    3
 5.05720229e-08-1.09413374e-11 4.82664708e+02 5.62014116e+01                   4
C6H5CH2OH               C   7H   8O   1     G    300.00   3500.00 1450.00      1
 1.25818433e+01 2.64134544e-02-7.93800081e-06 4.38368885e-10 8.64078241e-14    2
-1.87828960e+04-3.81332281e+01-6.02884966e+00 7.77532972e-02-6.10481830e-05    3
 2.48568434e-08-4.12367400e-12-1.33857950e+04 5.85676629e+01                   4
C6H5C2H                 C   8H   6          G    200.00   3500.00 1280.00      1
 1.52608075e+01 2.33328931e-02-9.12947266e-06 1.67060910e-09-1.19620465e-13    2
 3.14643486e+04-5.61979002e+01-2.98097335e+00 8.03384582e-02-7.59328693e-05    3
 3.64640448e-08-6.91521339e-12 3.61342445e+04 3.63113150e+01                   4
C6H4C2H                 C   8H   5          G    200.00   3500.00 1410.00      1
 1.60102851e+01 1.80276842e-02-6.10631304e-06 8.89485671e-10-4.39310966e-14    2
 6.01004864e+04-5.91795499e+01-2.59308035e+00 7.08031889e-02-6.22504670e-05    3
 2.74351849e-08-4.75061536e-12 6.53466354e+04 3.69628593e+01                   4
C6H5C2H3                C   8H   8          G    200.00   3500.00 1620.00      1
 2.08689866e+01 1.76153497e-02-4.02709770e-06 7.62327441e-11 4.96213672e-14    2
 7.92336643e+03-8.97908296e+01-4.75261300e+00 8.08785586e-02-6.26041430e-05    3
 2.41820127e-08-3.67040640e-12 1.62247647e+04 4.61791075e+01                   4
C6H5C2H5                C   8H  10          G    200.00   3500.00 1660.00      1
 2.15526198e+01 2.25377584e-02-5.71678900e-06 3.25230124e-10 3.67332240e-14    2
-7.08672334e+03-9.37205686e+01-4.75947959e+00 8.59404076e-02-6.30083395e-05    3
 2.33338849e-08-3.42842563e-12 1.64889366e+03 4.65555364e+01                   4
C6H5C2H2                C   8H   7          G    200.00   3500.00 1520.00      1
 1.92541492e+01 1.80154930e-02-5.00513538e-06 4.35360048e-10 9.55508855e-15    2
 3.83998805e+04-7.81182467e+01-4.29898223e+00 7.99974178e-02-6.61715085e-05    3
 2.72627167e-08-4.40283909e-12 4.55600324e+04 4.53739368e+01                   4
C6H5CHCH3               C   8H   9          G    200.00   3500.00 1700.00      1
 2.17404186e+01 1.87953835e-02-4.10980664e-06 2.52089055e-14 6.24670776e-14    2
 1.18126532e+04-9.21825542e+01-3.04486878e+00 7.71137068e-02-5.55671507e-05    3
 2.01793758e-08-2.90508448e-12 2.02396509e+04 4.05439039e+01                   4
XYLENE                  C   8H  10          G    200.00   3500.00 1800.00      1
 2.00142041e+01 2.37296538e-02-6.76483661e-06 7.09528579e-10-1.05910746e-14    2
-8.30085827e+03-8.55893397e+01-3.92128805e+00 7.69196362e-02-5.10898220e-05    3
 1.71261898e-08-2.29068292e-12 3.15918889e+02 4.39545368e+01                   4
RXYLENE                 C   8H   9          G    200.00   3500.00 1620.00      1
 2.04972472e+01 2.14206990e-02-5.61362499e-06 3.90127768e-10 2.53124037e-14    2
 1.19614473e+04-8.71674618e+01-3.85447681e+00 8.15484127e-02-6.12874339e-05    3
 2.33011602e-08-3.51034076e-12 1.98514059e+04 4.20634384e+01                   4
INDENE                  C   9H   8          G    200.00   3500.00 1610.00      1
 2.31048457e+01 1.91297559e-02-4.53547880e-06 1.22195972e-10 5.15079506e-14    2
 8.53092039e+03-1.04304485e+02-6.87762296e+00 9.36203612e-02-7.39366639e-05    3
 2.88597467e-08-4.41084465e-12 1.81852753e+04 5.46222710e+01                   4
INDENYL                 C   9H   7          G    200.00   3500.00 1430.00      1
 2.02650240e+01 2.20602663e-02-7.28401634e-06 9.93376351e-10-4.12200059e-14    2
 2.49669760e+04-8.59379510e+01-6.82385332e+00 9.78333498e-02-8.67662718e-05    3
 3.80480409e-08-6.51930821e-12 3.27143949e+04 5.44392226e+01                   4
C10H7                   C  10H   7          G    200.00   3500.00 1490.00      1
 2.12397133e+01 2.27484176e-02-6.96639984e-06 8.04033592e-10-1.68765509e-14    2
 3.76445828e+04-9.11799952e+01-6.45168846e+00 9.70877513e-02-8.18046553e-05    3
 3.42887116e-08-5.63511112e-12 4.58966205e+04 5.34576811e+01                   4
C10H7OH                 C  10H   8O   1     G    300.00   3500.00 1730.00      1
 2.61818201e+01 2.47079275e-02-8.75473292e-06 1.41213299e-09-8.61581287e-14    2
-1.58338679e+04-1.19314304e+02-3.09194587e+00 9.23929356e-02-6.74411561e-05    3
 2.40273250e-08-3.35424945e-12-5.70514485e+03 3.79602726e+01                   4
C10H7O                  C  10H   7O   1     G    200.00   3500.00 1520.00      1
 2.51245218e+01 2.12349548e-02-5.95579954e-06 5.14903131e-10 1.27934269e-14    2
 2.27944562e+03-1.11444322e+02-6.17635865e+00 1.03605693e-01-8.72427122e-05    3
 3.61670578e-08-5.85104780e-12 1.17949133e+04 5.26703345e+01                   4
C10H6CH3                C  11H   9          G    200.00   3500.00 1530.00      1
 2.52492992e+01 2.50352498e-02-6.91797983e-06 5.80759912e-10 1.70682319e-14    2
 3.22365783e+04-1.13732264e+02-6.94188380e+00 1.09195205e-01-8.94277403e-05    3
 3.65327252e-08-5.85743591e-12 4.20870803e+04 5.52614572e+01                   4
C10H7CH2                C  11H   9          G    200.00   3500.00 1480.00      1
 2.49658411e+01 2.73321300e-02-8.56499858e-06 1.05181162e-09-3.08780942e-14    2
 2.10853651e+04-1.11434380e+02-7.41870812e+00 1.14857939e-01-9.72735884e-05    3
 4.10106359e-08-6.78067949e-12 3.06711917e+04 5.74984562e+01                   4
C10H7CHO                C  11H   8O   1     G    200.00   3500.00 1700.00      1
 3.52801276e+01 1.31180777e-02-5.97592874e-07-9.89260930e-10 1.64133250e-13    2
-1.29136441e+04-1.70276966e+02-6.53399130e+00 1.11504240e-01-8.74089124e-05    3
 3.30543938e-08-4.84228656e-12 1.30315631e+03 5.36397397e+01                   4
C10H7CH3                C  11H  10          G    200.00   3500.00 1700.00      1
 3.19556728e+01 1.89589620e-02-2.92887011e-06-5.41540733e-10 1.30075404e-13    2
-1.51641367e+03-1.52538833e+02-7.17710562e+00 1.11036088e-01-8.41733928e-05    3
 3.13190564e-08-4.55530653e-12 1.17887310e+04 5.70191599e+01                   4
CH3C10H6OH              C  11H  10O   1     G    300.00   3500.00 1800.00      1
 2.91191897e+01 2.86451254e-02-9.80097852e-06 1.51373980e-09-8.72236902e-14    2
-2.13626722e+04-1.32660129e+02-1.76841840e+00 9.72842544e-02-6.70002527e-05    3
 2.26986562e-08-3.02957318e-12-1.02431333e+04 3.45100495e+01                   4
CH3C10H6O               C  11H   9O   1     G    300.00   3500.00 1800.00      1
 2.60936668e+01 3.24954890e-02-1.30480558e-05 2.52260734e-09-1.95492221e-13    2
-2.87397161e+03-1.14905163e+02-1.85059523e+00 9.45938490e-02-6.47966891e-05    3
 2.16887678e-08-2.85745896e-12 7.18596271e+03 3.63350123e+01                   4
C12H8                   C  12H   8          G    200.00   3500.00 1570.00      1
 2.77000844e+01 2.26169301e-02-5.57153301e-06 2.34722435e-10 5.00959715e-14    2
 1.79557617e+04-1.32407965e+02-8.95027502e+00 1.15993642e-01-9.47849520e-05    3
 3.81172783e-08-5.98215814e-12 2.94639745e+04 6.09409170e+01                   4
C12H7                   C  12H   7          G    200.00   3500.00 1550.00      1
 2.72643880e+01 2.07706230e-02-5.09002529e-06 1.94275307e-10 4.95145122e-14    2
 5.03500904e+04-1.28964283e+02-8.21375616e+00 1.12327124e-01-9.36930909e-05    3
 3.83031207e-08-6.09707346e-12 6.13483151e+04 5.77457264e+01                   4
BIPHENYL                C  12H  10          G    200.00   3500.00 1620.00      1
 3.03550359e+01 2.42378550e-02-5.78854421e-06 1.73422993e-10 6.27219799e-14    2
 7.33500793e+03-1.42781785e+02-7.48580998e+00 1.17672042e-01-9.23016807e-05    3
 3.57755368e-08-5.43143138e-12 1.95954420e+04 5.80338359e+01                   4
C12H9                   C  12H   9          G    300.00   3500.00 1430.00      1
 2.37129784e+01 3.27032248e-02-1.16108624e-05 1.80514888e-09-1.00355841e-13    2
 4.00500312e+04-1.02303917e+02-9.58279846e+00 1.25838265e-01-1.09304960e-04    3
 4.73501829e-08-8.06277438e-12 4.95726233e+04 7.02380080e+01                   4
FLUORENE                C  13H  10          G    200.00   3500.00 1580.00      1
 3.04982038e+01 2.54134231e-02-6.12248812e-06 2.13466649e-10 6.26037246e-14    2
 6.42405659e+03-1.44876977e+02-9.12300004e+00 1.25720268e-01-1.01350506e-04    3
 4.03940647e-08-6.29508585e-12 1.89443570e+04 6.43961517e+01                   4
C6H5CH2C6H5             C  13H  12          G    200.00   3500.00 1730.00      1
 3.68979008e+01 2.09448819e-02-2.15139957e-06-1.01983594e-09 1.90993633e-13    2
 1.61235186e+03-1.77722084e+02-9.21937277e+00 1.27574416e-01-9.46047530e-05    3
 3.46076605e-08-4.95748852e-12 1.75689285e+04 7.00449671e+01                   4
C14H10                  C  14H  10          G    200.00   3500.00 1550.00      1
 3.33910437e+01 2.79675435e-02-7.16204131e-06 3.82999815e-10 5.29487368e-14    2
 8.53645744e+03-1.60739802e+02-9.79770432e+00 1.39422377e-01-1.15021558e-04    3
 4.67741896e-08-7.42950123e-12 2.19249693e+04 6.65486230e+01                   4
C14H9                   C  14H   9          G    298.15   3500.00 1380.00      1
 2.51054798e+01 4.12375740e-02-1.71094085e-05 3.35330087e-09-2.55891930e-13    2
 4.20489547e+04-1.12231126e+02-1.15966330e+01 1.47620510e-01-1.32743034e-04    3
 5.92149558e-08-1.03757570e-11 5.21787378e+04 7.66564973e+01                   4
C16H10                  C  16H  10          G    200.00   3500.00 1560.00      1
 3.81807384e+01 2.83119132e-02-6.73304717e-06 1.57163103e-10 8.21180996e-14    2
 9.09208783e+03-1.88517734e+02-1.17161987e+01 1.56252778e-01-1.29753109e-04    3
 5.27298391e-08-8.34299024e-12 2.46599322e+04 7.43946050e+01                   4
C16H9                   C  16H   9          G    300.00   3500.00 1240.00      1
 1.61933943e+01 6.96117237e-02-3.71054209e-05 9.43826309e-09-9.32516221e-13    2
 4.61008367e+04-6.54256061e+01-1.33382682e+01 1.64875151e-01-1.52343438e-04    3
 7.13941862e-08-1.34236298e-11 5.34246890e+04 8.34001912e+01                   4
C6H5C2H4C6H5            C  14H  14          G    300.00   3500.00 1170.00      1
 6.79293376e+00 9.36089877e-02-5.25184338e-05 1.38852177e-08-1.40951786e-12    2
 1.04787081e+04-8.65156409e+00-1.16088783e+01 1.56521166e-01-1.33175072e-04    3
 5.98434163e-08-1.12296458e-11 1.47847321e+04 8.30156954e+01                   4
C18H10                  C  18H  10          G    300.00   3500.00 1430.00      1
 3.55205983e+01 2.97059186e-02-5.18577074e-06-7.74977698e-10 2.05764425e-13    2
 1.13998029e+04-1.72584660e+02-1.43149515e+01 1.69106058e-01-1.51409693e-04    3
 6.73946831e-08-1.17120084e-11 2.56527702e+04 8.56679626e+01                   4
C18H9                   C  18H   9          G    300.00   3500.00 1110.00      1
 1.00826785e+01 9.26185724e-02-5.34378503e-05 1.44603230e-08-1.49786384e-12    2
 4.90427509e+04-3.41228910e+01-1.54340435e+01 1.84570724e-01-1.77697514e-04    3
 8.90907519e-08-1.83065190e-11 5.47074632e+04 9.16434681e+01                   4
LC6H5                   C   6H   5          G    300.00   3500.00 1140.00      1
 1.23076079e+01 1.68261942e-02-6.51181276e-06 1.21158858e-09-8.99427818e-14    2
 5.89425071e+04-3.55373263e+01 1.67614201e-01 5.94226632e-02-6.25597982e-05    3
 3.39881883e-08-7.27779359e-12 6.17104257e+04 2.46218078e+01                   4
C6H2                    C   6H   2          G    200.00   3500.00  700.00      1
 9.95239950e+00 1.43744769e-02-7.32585513e-06 1.80931756e-09-1.74471724e-13    2
 8.06473021e+04-2.49945451e+01-5.39476048e-01 7.43280514e-02-1.35797801e-04    3
 1.24163551e-07-4.38724124e-11 8.21161647e+04 2.18805005e+01                   4
C6H3                    C   6H   3          G    300.00   3500.00 1320.00      1
 1.19194526e+01 1.16137824e-02-4.19264458e-06 6.84692858e-10-4.17887320e-14    2
 8.26280759e+04-3.29876558e+01 4.46601449e+00 3.41999584e-02-2.98587536e-05    3
 1.36473742e-08-2.49684202e-12 8.45957836e+04 5.04018540e+00                   4
C6H4                    C   6H   4          G    300.00   3500.00 1360.00      1
 1.74447671e+01 6.21306801e-03-9.80964592e-07 8.00596955e-11-2.88323342e-15    2
 5.49568895e+04-6.59208062e+01-1.17305602e+00 6.09713714e-02-6.13761521e-05    3
 2.96855438e-08-5.44506781e-12 6.00209374e+04 2.96241241e+01                   4
C8H2                    C   8H   2          G    300.00   3500.00 1060.00      1
 1.62719352e+01 9.99874486e-03-2.93037073e-06 2.89537311e-10 2.52409677e-16    2
 1.07885459e+05-5.89733616e+01 1.87361702e-01 7.06952486e-02-8.88216496e-05    3
 5.43092096e-08-1.27402363e-11 1.11295389e+05 1.95626383e+01                   4
BIN1B                   C  20H  10          G    300.00   3500.00 1430.00      1
 3.76362472e+01 4.45434591e-02-1.43416639e-05 1.85353170e-09-6.45806827e-14    2
-9.82259049e+02-1.87789152e+02-1.59101511e+01 1.94323594e-01-1.71453694e-04    3
 7.50992333e-08-1.28697733e-11 1.43320109e+04 8.96934452e+01                   4
BIN1A                   C  20H  16          G    300.00   3500.00 1410.00      1
 4.18190040e+01 5.54173380e-02-1.89314361e-05 2.76164477e-09-1.34640474e-13    2
-3.16800626e+03-2.10125772e+02-1.45702447e+01 2.15386838e-01-1.89111755e-04    3
 8.32251525e-08-1.44012199e-11 1.27337619e+04 8.12945223e+01                   4
C18H14                  H  14C  18          G    100.00   3500.00  700.00      1
-8.78909820e+00 1.54177573e-01-9.84392856e-05 2.89551421e-08-3.12416384e-12    2
 3.49494076e+04 6.52592559e+01-7.00582258e+00 1.43987427e-01-7.66032577e-05    3
 8.15892501e-09 4.30305656e-12 3.46997490e+04 5.72920316e+01                   4
C6H5C2H4                C   8H   9          G    200.00   3500.00 1530.00      1
 1.90733225e+01 2.32393266e-02-7.04814960e-06 8.06137047e-10-1.68210968e-14    2
 1.95612169e+04-7.66267073e+01-3.58296935e+00 8.24714621e-02-6.51188707e-05    3
 2.61092835e-08-4.15132215e-12 2.64940422e+04 4.23117942e+01                   4
RMCYC6                  C   7H  13          G    300.00   3500.00 1800.00      1
 1.73339089e+01 3.85260766e-02-1.58310783e-05 3.15191350e-09-2.53163676e-13    2
-5.89958084e+03-7.33836570e+01-9.95790350e+00 9.91745487e-02-6.63714717e-05    3
 2.18705777e-08-2.85297815e-12 3.92547164e+03 7.43253253e+01                   4
MCYC6                   C   7H  14          G    300.00   3500.00 1800.00      1
 1.67194642e+01 4.36180495e-02-1.87773262e-05 3.92058734e-09-3.26702691e-13    2
-2.91866329e+04-7.40612288e+01-1.01006365e+01 1.03218273e-01-6.84441793e-05    3
 2.23157181e-08-2.88158197e-12-1.95313966e+04 7.10947511e+01                   4
TMBENZ                  C   9H  12          G    300.00   3500.00 1800.00      1
 1.47576863e+01 4.50315820e-02-1.97554191e-05 4.21197805e-09-3.57314904e-13    2
-1.09025840e+04-5.35378410e+01-2.75522788e+00 8.39491691e-02-5.21867417e-05    3
 1.62235790e-08-2.02559281e-12-4.59793488e+03 4.12457040e+01                   4
NPBENZ                  C   9H  12          G    300.00   3500.00 1600.00      1
 1.88963385e+01 3.80090263e-02-1.52789365e-05 2.95630025e-09-2.27699137e-13    2
-8.96605333e+03-7.62711351e+01-5.58650169e+00 9.92161268e-02-7.26605932e-05    3
 2.68653239e-08-3.96348408e-12-1.13154446e+03 5.33514402e+01                   4
RC9H11                  C   9H  11          G    300.00   3500.00 1800.00      1
 1.94777753e+01 3.52558754e-02-1.42493119e-05 2.76058036e-09-2.13044853e-13    2
 6.10938509e+03-7.94714191e+01-1.83523076e+00 8.26181111e-02-5.37178417e-05    3
 1.73785543e-08-2.24331902e-12 1.37820673e+04 3.58790159e+01                   4
DIBZFUR                 C  12H   8O   1     G    300.00   3500.00 1410.00      1
 2.49525253e+01 3.24730740e-02-1.15459384e-05 1.79679089e-09-9.97834068e-14    2
-5.30753643e+03-1.13355891e+02-1.16970901e+01 1.36443614e-01-1.22152896e-04    3
 5.40932247e-08-9.37220075e-12 5.02765511e+03 7.60497479e+01                   4
BZFUR                   C   8H   6O   1     G    300.00   3500.00 1380.00      1
 1.64578320e+01 2.37623599e-02-8.52218857e-06 1.36123792e-09-7.97160791e-14    2
-5.90596930e+03-6.59480309e+01-8.70136925e+00 9.66875810e-02-8.77887332e-05    3
 3.96542547e-08-7.01685679e-12 1.03797025e+03 6.35339354e+01                   4
ODECAL                  C  10H  18          G    300.00   3500.00 1800.00      1
 2.82109951e+01 4.74108378e-02-1.82963840e-05 3.42084129e-09-2.57817094e-13    2
-2.68355233e+04-1.31410209e+02-1.02710770e+01 1.32926554e-01-8.95594805e-05    3
 2.98145807e-08-3.92361424e-12-1.29819774e+04 7.68627935e+01                   4
DECALIN                 C  10H  18          G    300.00   3500.00 1750.00      1
 2.70110184e+01 4.68748410e-02-1.63895662e-05 2.62564196e-09-1.59790271e-13    2
-3.79226248e+04-1.35167686e+02-1.45870776e+01 1.41956203e-01-9.78878768e-05    3
 3.36726175e-08-4.59507248e-12-2.33632912e+04 8.87980329e+01                   4
TETRALIN                C  10H  12          G    300.00   3500.00 1650.00      1
 2.40250650e+01 3.45031755e-02-1.26565584e-05 2.20632612e-09-1.51941366e-13    2
-9.85314234e+03-1.11161754e+02-1.00807334e+01 1.17183899e-01-8.78208525e-05    3
 3.25757379e-08-4.75336739e-12 1.40177115e+03 7.04583491e+01                   4
DCYC5                   C  10H  16          G    300.00   3500.00 1750.00      1
 2.70110184e+01 4.68748410e-02-1.63895662e-05 2.62564196e-09-1.59790271e-13    2
-3.79226248e+04-1.35167686e+02-1.45870776e+01 1.41956203e-01-9.78878768e-05    3
 3.36726175e-08-4.59507248e-12-2.33632912e+04 8.87980329e+01                   4
RTETRALIN               C  10H  11          G    300.00   3500.00 1800.00      1
 2.92427993e+01 2.67836077e-02-9.17250453e-06 1.42952815e-09-8.46469052e-14    2
 3.95646759e+03-1.44540573e+02-1.09331570e+01 1.16063511e-01-8.35724236e-05    3
 2.89850537e-08-3.91180323e-12 1.84198119e+04 7.29000838e+01                   4
RTETRAOO                C  10H  11O   2     G    300.00   3500.00 1800.00      1
 5.34619204e+01-7.89286507e-03 1.09697433e-05-3.89490463e-09 4.38586931e-13    2
-1.76924226e+04-2.71823519e+02-1.36343940e+01 1.41210056e-01-1.13282691e-04    3
 4.21245154e-08-5.95299919e-12 6.46225063e+03 9.13157320e+01                   4
RDECALIN                C  10H  17          G    300.00   3500.00 1800.00      1
 2.85620385e+01 4.11366283e-02-1.36024033e-05 2.01592555e-09-1.09376388e-13    2
-1.53025082e+04-1.39641715e+02-1.39601311e+01 1.35630338e-01-9.23471617e-05    3
 3.11806509e-08-4.16003269e-12 5.47280143e+00 9.04971374e+01                   4
RODECA                  C  10H  17          G    300.00   3500.00 1800.00      1
 2.85620385e+01 4.11366283e-02-1.36024033e-05 2.01592555e-09-1.09376388e-13    2
-1.53025082e+04-1.39641715e+02-1.39601311e+01 1.35630338e-01-9.23471617e-05    3
 3.11806509e-08-4.16003269e-12 5.47280143e+00 9.04971374e+01                   4
NC10H22                 C  10H  22          G    300.00   3500.00 1800.00      1
 2.92878820e+01 5.29921188e-02-1.98404688e-05 3.55616754e-09-2.54281575e-13    2
-4.56232341e+04-1.22751993e+02-2.17870059e+00 1.22917858e-01-7.81119181e-05    3
 2.51381858e-08-3.25178411e-12-3.42952644e+04 4.75517162e+01                   4
NC10H21                 C  10H  21          G    300.00   3500.00 1800.00      1
 2.63212767e+01 5.52219590e-02-2.21266426e-05 4.33498609e-09-3.42316219e-13    2
-2.10175200e+04-1.03193018e+02-1.81057340e+00 1.17737181e-01-7.42226612e-05    3
 2.36298078e-08-3.02215257e-12-1.08900539e+04 4.90624235e+01                   4
C10H10                  C  10H  10          G    300.00   3500.00 1800.00      1
 1.82592674e+01 4.15934266e-02-1.83631866e-05 3.88491233e-09-3.27420909e-13    2
 4.39687909e+03-8.23923085e+01-1.14588962e+01 1.07633790e-01-7.33968229e-05    3
 2.42677406e-08-3.15836928e-12 1.50954180e+04 7.84485924e+01                   4
NC12H25                 C  12H  25          G    300.00   3500.00 1800.00      1
 3.17005400e+01 6.61544689e-02-2.66295479e-05 5.21805220e-09-4.10999243e-13    2
-2.88525830e+04-1.31607526e+02-2.06085002e+00 1.41179780e-01-8.91506405e-05    3
 2.83740124e-08-3.62710483e-12-1.66984826e+04 5.11161596e+01                   4
IC16H33                 C  16H  33          G    300.00   3500.00 1650.00      1
 5.11453797e+01 7.53296293e-02-2.79262920e-05 4.92907249e-09-3.44363400e-13    2
-5.61938948e+04-2.43048347e+02-8.95216391e+00 2.21020644e-01-1.60372669e-04    3
 5.84427602e-08-8.45249790e-12-3.63617054e+04 7.69829261e+01                   4
NC16H33                 C  16H  33          G    300.00   3500.00 1800.00      1
 4.66278463e+01 8.00212049e-02-3.03236203e-05 5.55903238e-09-4.09822165e-13    2
-4.61545245e+04-2.04019531e+02-3.22413441e+00 1.90803384e-01-1.22642103e-04    3
 3.97510631e-08-5.15871531e-12-2.82078114e+04 6.57897888e+01                   4
NC10H19                 C  10H  19          G    300.00   3500.00 1800.00      1
 9.88286994e+00 2.86275431e-02-1.23662483e-05 2.58308667e-09-2.14521125e-13    2
 7.14211786e+03-2.81379541e+01-9.61360365e-01 5.27258326e-02-3.24481563e-05    3
 1.00208304e-08-1.24754108e-12 1.10460408e+04 3.05532826e+01                   4
NC12H26                 C  12H  26          G    300.00   3500.00 1800.00      1
 3.61414017e+01 6.11046044e-02-2.24641185e-05 3.93182761e-09-2.73349693e-13    2
-5.40359156e+04-1.56831918e+02-2.66627653e+00 1.47343889e-01-9.43301893e-05    3
 3.05488909e-08-3.97016404e-12-4.00651514e+04 5.32033327e+01                   4
IC16H34                 C  16H  34          G    300.00   3500.00 1590.00      1
 4.72524577e+01 8.54680800e-02-3.36612750e-05 6.38202103e-09-4.82094960e-13    2
-7.78744134e+04-2.24182938e+02-9.93612209e+00 2.29338721e-01-1.69388295e-04    3
 6.32906247e-08-9.42998862e-12-5.96884450e+04 7.82391913e+01                   4
NC16H34                 C  16H  34          G    300.00   3500.00 1800.00      1
 4.98210209e+01 7.73881742e-02-2.77557933e-05 4.69678208e-09-3.12959347e-13    2
-7.08514653e+04-2.24842840e+02-3.64057950e+00 1.96191731e-01-1.26758757e-04    3
 4.13645464e-08-5.40570439e-12-5.16052891e+04 6.45024943e+01                   4
NC10H20                 C  10H  20          G    300.00   3500.00 1800.00      1
 2.82971765e+01 4.89478994e-02-1.82737102e-05 3.23575318e-09-2.26811965e-13    2
-3.12534572e+04-1.16784043e+02-2.31417696e+00 1.16973129e-01-7.49614017e-05    3
 2.42311945e-08-3.14284548e-12-2.02333700e+04 4.88909872e+01                   4
IC12H26                 C  12H  26          G    300.00   3500.00 1800.00      1
 3.61414017e+01 6.11046044e-02-2.24641185e-05 3.93182761e-09-2.73349693e-13    2
-5.40359156e+04-1.56831918e+02-2.66627653e+00 1.47343889e-01-9.43301893e-05    3
 3.05488909e-08-3.97016404e-12-4.00651514e+04 5.32033327e+01                   4
IC12H25                 C  12H  25          G    300.00   3500.00 1800.00      1
 3.17005400e+01 6.61544689e-02-2.66295479e-05 5.21805220e-09-4.10999243e-13    2
-2.88525830e+04-1.31607526e+02-2.06085002e+00 1.41179780e-01-8.91506405e-05    3
 2.83740124e-08-3.62710483e-12-1.66984826e+04 5.11161596e+01                   4
C10H16                  C  10H  16          G    300.00   3500.00 1800.00      1
 2.89286842e+01 4.33698796e-02-1.66040875e-05 3.00058304e-09-2.14827238e-13    2
-2.62353997e+04-1.44986797e+02-1.64117642e+01 1.44126432e-01-1.00567881e-04    3
 3.40982842e-08-4.53395241e-12-9.91283830e+03 1.00405168e+02                   4
C10H15                  C  10H  15          G    300.00   3500.00 1770.00      1
 3.20501518e+01 3.53882668e-02-1.22004910e-05 1.87186805e-09-1.05121849e-13    2
-9.38258806e+03-1.63611813e+02-1.67888466e+01 1.45758885e-01-1.05734913e-04    3
 3.71014055e-08-5.08104522e-12 7.90641738e+03 9.98941922e+01                   4
C6H5C4H9                C  10H  14          G    300.00   3500.00 1620.00      1
 2.20508185e+01 4.25105669e-02-1.68597803e-05 3.21475888e-09-2.44036189e-13    2
-1.30455889e+04-9.17624124e+01-5.81141693e+00 1.11306210e-01-8.05594497e-05    3
 2.94286146e-08-4.28938429e-12-4.01822460e+03 5.60982384e+01                   4
RC6H5C4H8               C  10H  13          G    300.00   3500.00 1650.00      1
 2.28150931e+01 3.94891629e-02-1.56943246e-05 2.97948476e-09-2.24328474e-13    2
 4.22312781e+03-9.69374998e+01-3.49464093e+00 1.03270336e-01-7.36772096e-05    3
 2.64069130e-08-3.77393882e-12 1.29053401e+04 4.31670233e+01                   4
C6H5C4H7-3              C  10H  12          G    300.00   3500.00 1480.00      1
 1.62604487e+01 4.74926281e-02-2.11208381e-05 4.52916148e-09-3.83728373e-13    2
 2.53220514e+03-5.97389803e+01-5.26848528e+00 1.05678936e-01-8.00934476e-05    3
 3.10934000e-08-4.87093083e-12 8.90476960e+03 5.25659295e+01                   4
CH2OHCH2OH              C   2H   6O   2     G    300.00   3500.00 1510.00      1
 8.58229296e+00 1.47365723e-02-4.87454239e-06 7.03407917e-10-3.54291327e-14    2
-5.09140292e+04-1.61663174e+01-4.19778996e-01 3.85831205e-02-2.85631665e-05    3
 1.11619616e-08-1.76697775e-12-4.81954035e+04 3.09733168e+01                   4
GLYCEROL                C   3H   8O   3     G    300.00   3500.00 1260.00      1
 1.38765800e+01 2.06689875e-02-7.56631316e-06 1.26540543e-09-8.07917221e-14    2
-7.51651917e+04-3.83652390e+01 3.56065367e+00 5.34179599e-02-4.65531851e-05    3
 2.18933800e-08-4.17364382e-12-7.25655783e+04 1.37872737e+01                   4
C3H4O3                  C   3H   4O   3     G    300.00   3500.00 1710.00      1
 1.37242814e+01 1.08811102e-02-3.70124803e-06 5.78901295e-10-3.43205672e-14    2
-5.77802808e+04-3.99570095e+01 2.17563099e+00 3.78954972e-02-2.73980787e-05    3
 9.81743178e-09-1.38498292e-12-5.38306424e+04 2.19543276e+01                   4
FURFURAL                C   5H   4O   2     G    300.00   3500.00 1430.00      1
 1.05158973e+01 2.23224204e-02-1.09267077e-05 2.56683180e-09-2.34844936e-13    2
-2.33303223e+04-2.94000431e+01-1.81996663e+00 5.68283336e-02-4.71217216e-05    3
 1.94409641e-08-3.18486807e-12-1.98022652e+04 3.45255930e+01                   4
FURAN                   C   4H   4O   1     G    300.00   3500.00 1250.00      1
 8.37486474e+00 1.95634449e-02-9.90167102e-06 2.37694376e-09-2.20517691e-13    2
-9.41817582e+03-2.52053388e+01-7.59507782e+00 7.06672610e-02-7.12262504e-05    3
 3.50833861e-08-6.76180616e-12-5.42569018e+03 5.54039922e+01                   4
CH2CCHCHO               C   4H   4O   1     G    300.00   3500.00 1590.00      1
 1.05858587e+01 1.29955935e-02-4.76360657e-06 7.49448020e-10-3.96845891e-14    2
 3.10513221e+03-2.93262571e+01 1.05971995e+00 3.69607224e-02-2.73722187e-05    3
 1.02289500e-08-1.53017232e-12 6.13444432e+03 2.10494502e+01                   4
C4H3O                   C   4H   3O   1     G    300.00   3500.00 1240.00      1
 8.44125951e+00 1.62911123e-02-8.34126337e-06 2.01436734e-09-1.87394567e-13    2
 1.94535774e+04-2.27855102e+01-5.90872261e+00 6.25813772e-02-6.43375516e-05    3
 3.21198986e-08-6.25705813e-12 2.30123730e+04 4.95317029e+01                   4
MEFU2                   C   5H   6O   1     G    300.00   3500.00 1260.00      1
 5.16398130e+00 3.29529092e-02-1.68209206e-05 4.03716089e-09-3.55511413e-13    2
-1.31841669e+04-2.67616512e+00-3.74149807e+00 6.12242723e-02-5.04773052e-05    3
 2.18447718e-08-3.88876755e-12-1.09399861e+04 4.23457857e+01                   4
DMF                     C   6H   8O   1     G    300.00   3500.00 1590.00      1
 1.38889512e+01 2.49736910e-02-8.98420928e-06 1.42738209e-09-7.97717653e-14    2
-2.20872036e+04-4.94041143e+01-2.31533190e+00 6.57391831e-02-4.74422206e-05    3
 1.75523344e-08-2.61514163e-12-1.69342416e+04 3.62866619e+01                   4
DMF-3YL                 C   6H   7O   1     G    300.00   3500.00 1620.00      1
 1.41703390e+01 2.18230103e-02-7.69511491e-06 1.17891326e-09-6.12376920e-14    2
 1.19557794e+04-4.86583466e+01-1.12307983e+00 5.95845384e-02-4.26594928e-05    3
 1.55675461e-08-2.28170573e-12 1.69108471e+04 3.25015042e+01                   4
C6H10O5                 C   6H  10O   5     G    300.00   3500.00 1220.00      1
 1.54889701e+01 4.96354436e-02-2.45944552e-05 5.82332728e-09-5.35666028e-13    2
-1.09180509e+05-4.81819746e+01-7.95116443e+00 1.26488344e-01-1.19085726e-04    3
 5.74579013e-08-1.11165214e-11-1.03461116e+05 6.95642156e+01                   4
C6H8O4                  C   6H   8O   4     G    300.00   3500.00 1300.00      1
 1.58073737e+01 3.77998802e-02-1.77241244e-05 3.97559911e-09-3.49009601e-13    2
-7.78788475e+04-5.15128466e+01-4.55493859e+00 1.00453149e-01-9.00163573e-05    3
 4.10485391e-08-7.47842113e-12-7.25846463e+04 5.20658826e+01                   4
C6H6O3                  C   6H   6O   3     G    300.00   3500.00 1770.00      1
 1.98638064e+01 1.79335036e-02-5.95409002e-06 8.93594360e-10-4.95460319e-14    2
-4.95264841e+04-7.44496641e+01 7.10718650e-01 6.12173177e-02-4.26352883e-05    3
 1.47094883e-08-2.00094348e-12-4.27462910e+04 2.88889339e+01                   4
C5H8O4                  C   5H   8O   4     G    300.00   3500.00 1230.00      1
 1.19601516e+01 3.99450904e-02-1.95947427e-05 4.60940299e-09-4.22302501e-13    2
-8.26385853e+04-2.91875110e+01-6.95683226e+00 1.01463737e-01-9.46174827e-05    3
 4.52721347e-08-8.68708537e-12-7.79850073e+04 6.59920850e+01                   4
CATECHOL                C   6H   6O   2     G    300.00   3500.00 1150.00      1
 1.43499786e+01 2.44086069e-02-1.04210986e-05 2.01939014e-09-1.47232869e-13    2
-3.94515396e+04-4.76262801e+01-5.49815252e+00 9.34455847e-02-1.00469330e-04    3
 5.42212637e-08-1.14954663e-11-3.48864694e+04 5.09034926e+01                   4
GUAIACOL                C   7H   8O   2     G    300.00   3500.00 1000.00      1
 9.99301768e+00 4.50609487e-02-2.36180832e-05 5.74985949e-09-5.33615067e-13    2
-3.55531887e+04-2.30989126e+01-7.52910606e+00 1.15149444e-01-1.28750826e-04    3
 7.58383544e-08-1.80557388e-11-3.20487639e+04 6.14352057e+01                   4
SALICALD                C   7H   6O   2     G    300.00   3500.00 1580.00      1
 2.23242879e+01 1.54051217e-02-2.83991362e-06-4.41656070e-10 1.22876830e-13    2
-3.64536806e+04-8.95534716e+01-5.00623414e+00 8.45963168e-02-6.85277571e-05    3
 2.72747336e-08-4.26262786e-12-2.78172356e+04 5.48021588e+01                   4
VANILLIN                C   8H   8O   3     G    300.00   3500.00 1260.00      1
 1.36544659e+01 4.84143197e-02-2.42641766e-05 5.50487717e-09-4.76001813e-13    2
-5.18855419e+04-3.54575775e+01-4.86637432e+00 1.07210638e-01-9.42597935e-05    3
 4.25395951e-08-7.82416013e-12-4.72182901e+04 5.81751538e+01                   4
C8H6O3                  C   8H   6O   3     G    300.00   3500.00 1000.00      1
 4.59309000e+00 6.23299032e-02-3.47374634e-05 8.74937443e-09-8.39789258e-13    2
-4.48191761e+04 1.51136238e+01-8.47052147e+00 1.14584349e-01-1.13119132e-04    3
 6.10038203e-08-1.39034007e-11-4.22064538e+04 7.81379977e+01                   4
C6H5OCH3                C   7H   8O   1     G    300.00   3500.00 1380.00      1
 1.25085131e+01 3.49906136e-02-1.63096094e-05 3.64836870e-09-3.19988435e-13    2
-1.52038793e+04-4.20406469e+01-5.29461544e+00 8.65938847e-02-7.24001214e-05    3
 3.07452344e-08-5.22884092e-12-1.02902158e+04 4.95832509e+01                   4
C7H6O3                  C   7H   6O   3     G    300.00   3500.00 1000.00      1
 9.61003547e+00 4.63126478e-02-2.49854435e-05 6.23130958e-09-5.96781904e-13    2
-5.28813089e+04-1.46625797e+01-7.07010612e+00 1.13033214e-01-1.25066293e-04    3
 7.29518760e-08-1.72769235e-11-4.95452806e+04 6.58094615e+01                   4
RC7H5O3                 C   7H   5O   3     G    300.00   3500.00 1000.00      1
 1.03519979e+01 4.06949748e-02-2.16398118e-05 5.16863274e-09-4.69580354e-13    2
-3.48541025e+04-1.78724726e+01-6.94106362e+00 1.09867221e-01-1.25398181e-04    3
 7.43408789e-08-1.77626419e-11-3.13954902e+04 6.55565530e+01                   4
C24H28O4                C  24H  28O   4     G    300.00   3500.00 1080.00      1
 1.29252082e+01 8.11297206e-02-4.64957344e-05 1.23575596e-08-1.22239418e-12    2
-7.66058398e+03-2.94388861e+00 3.08710559e+00 1.17567138e-01-9.71032581e-05    3
 4.35967718e-08-8.45369329e-12-5.53555382e+03 4.52764201e+01                   4
C6H4O                   C   6H   4O   1     G    300.00   3500.00 1320.00      1
 1.34428169e+01 1.79658727e-02-6.67332756e-06 1.12237508e-09-7.10809389e-14    2
 1.54076839e+04-4.72500521e+01-4.80707073e+00 7.32685624e-02-6.95172932e-05    3
 3.28617516e-08-6.08232650e-12 2.02256542e+04 4.58618541e+01                   4
RSALICPH                C   7H   5O   2     G    300.00   3500.00 1000.00      1
 6.00653602e+00 4.55336022e-02-2.51852434e-05 6.39158447e-09-6.19568333e-13    2
 4.68000652e+02 2.82366759e+00-8.00629333e+00 1.01584920e-01-1.09262219e-04    3
 6.24429019e-08-1.46323977e-11 3.27056652e+03 7.04274690e+01                   4
RGUAIPH                 C   7H   7O   2     G    300.00   3500.00 1000.00      1
 1.03288611e+01 4.15815421e-02-2.20221217e-05 5.39151141e-09-5.01575158e-13    2
-4.91455292e+03-2.20047788e+01-7.23884843e+00 1.11852380e-01-1.27428379e-04    3
 7.56623495e-08-1.80692847e-11-1.40101102e+03 6.27492646e+01                   4
RANISPH                 C   7H   7O   1     G    300.00   3500.00 1000.00      1
 6.14038303e+00 4.52741710e-02-2.46495251e-05 6.30633051e-09-6.15603088e-13    2
 1.78813934e+04-4.35386479e+00-8.02841886e+00 1.01949379e-01-1.09662336e-04    3
 6.29815381e-08-1.47844050e-11 2.07151538e+04 6.40024140e+01                   4
RCATEPH                 C   6H   5O   2     G    300.00   3500.00 1000.00      1
 1.18218903e+01 2.70911140e-02-1.34162461e-05 3.08575127e-09-2.72412036e-13    2
-7.82412444e+03-3.10506037e+01-7.41421142e+00 1.04035521e-01-1.28832857e-04    3
 8.00301583e-08-1.95085138e-11-3.97690409e+03 6.17524678e+01                   4
CH3OCH3                 C   2H   6O   1     G    300.00   3500.00 1800.00      1
 4.75053937e+00 1.85969231e-02-7.67398928e-06 1.52676702e-09-1.21721527e-13    2
-2.48946039e+04-1.32907051e+00 8.26271820e-01 2.73175177e-02-1.49411514e-05    3
 4.21830855e-09-4.95546740e-13-2.34818676e+04 1.99098841e+01                   4
CH3OCH2                 C   2H   5O   1     G    300.00   3500.00 1800.00      1
 4.38698121e+00 1.62462160e-02-6.72869512e-06 1.35709467e-09-1.09478883e-13    2
-2.38681615e+03 3.59289931e+00 1.56125465e+00 2.25256083e-02-1.19615221e-05    3
 3.29517873e-09-3.78657225e-13-1.36955459e+03 1.88863209e+01                   4
DME-OO                  C   2H   5O   3     G    300.00   3500.00 1800.00      1
 1.28946522e+01 1.03828333e-02-3.02554925e-06 3.64876465e-10-1.24114560e-14    2
-2.39005723e+04-3.76069422e+01 3.24067850e+00 3.18361082e-02-2.09032783e-05    3
 6.98625761e-09-9.32047726e-13-2.04251417e+04 1.46423774e+01                   4
DME-QOOH                C   2H   5O   3     G    300.00   3500.00 1250.00      1
 1.07374986e+01 1.39769737e-02-5.32012511e-06 9.94916291e-10-7.50060773e-14    2
-1.73025110e+04-2.35990452e+01 1.12063957e-01 4.79783647e-02-4.61217943e-05    3
 2.27558065e-08-4.42718413e-12-1.46461523e+04 3.00335324e+01                   4
DME-OOQOOH              C   2H   5O   5     G    300.00   3500.00 1370.00      1
 1.59411134e+01 1.44932658e-02-5.65696988e-06 1.09027769e-09-8.49010010e-14    2
-3.74943653e+04-4.65328770e+01 2.39014292e+00 5.40581429e-02-4.89761785e-05    3
 2.21701845e-08-3.93159933e-12-3.37813994e+04 2.31087131e+01                   4
DME-OQOOH               C   2H   4O   4     G    300.00   3500.00 1760.00      1
 1.54960902e+01 1.58757331e-03 2.24426442e-06-9.74238763e-10 1.03773225e-13    2
-4.69655446e+04-5.18401371e+01 3.62388925e+00 2.85698483e-02-2.07519927e-05    3
 7.73646468e-09-1.13354260e-12-4.27865299e+04 1.21478891e+01                   4
MTBE                    C   5H  12O   1     G    300.00   3500.00 1320.00      1
 9.85250850e+00 4.01896196e-02-1.66704212e-05 3.10158953e-09-2.11537800e-13    2
-4.09274217e+04-2.61941107e+01-1.85856421e+00 7.56777187e-02-5.69978066e-05    3
 2.34689559e-08-4.06899355e-12-3.78356985e+04 3.35564109e+01                   4
ETBE                    C   6H  14O   1     G    300.00   3500.00 1280.00      1
 1.16559129e+01 4.67934007e-02-1.93342030e-05 3.59185193e-09-2.45565035e-13    2
-4.60322111e+04-3.38084898e+01-3.48005590e+00 9.40933031e-02-7.47637761e-05    3
 3.24614212e-08-5.88415279e-12-4.21574031e+04 4.29502764e+01                   4
DIPE                    C   6H  14O   1     G    300.00   3500.00 1380.00      1
 1.11573938e+01 4.99175632e-02-2.25561365e-05 4.38444774e-09-3.06549287e-13    2
-4.59357932e+04-3.06117818e+01-2.50745285e+00 8.95258145e-02-6.56085835e-05    3
 2.51827313e-08-4.07435429e-12-4.21642955e+04 3.97144261e+01                   4
TAME                    C   6H  14O   1     G    300.00   3500.00 1320.00      1
 1.13309755e+01 4.74280959e-02-1.96957514e-05 3.66860789e-09-2.50688272e-13    2
-4.42745213e+04-3.17952363e+01-2.12836714e+00 8.82139827e-02-6.60433501e-05    3
 2.70764860e-08-4.68399852e-12-4.07212548e+04 3.68750524e+01                   4
RMTBE                   C   5H  11O   1     G    300.00   3500.00 1370.00      1
 1.09269218e+01 3.74766294e-02-1.73062498e-05 3.86241491e-09-3.39119828e-13    2
-1.88007824e+04-2.53563622e+01-1.81069336e-01 6.99087204e-02-5.28158384e-05    3
 2.11420201e-08-3.49233245e-12-1.57571928e+04 3.17301890e+01                   4
RDIPE                   C   6H  13O   1     G    300.00   3500.00 1800.00      1
 1.69549485e+01 3.45118442e-02-1.31342745e-05 2.36150251e-09-1.67133165e-13    2
-2.78147474e+04-5.54607929e+01 6.91787229e-01 7.06522026e-02-4.32512399e-05    3
 1.35159341e-08-1.71635978e-12-2.19600093e+04 3.25588286e+01                   4
MTBE-O                  C   5H  10O   2     G    300.00   3500.00 1520.00      1
 1.51388761e+01 2.99979376e-02-1.22799221e-05 2.46100792e-09-1.97690787e-13    2
-5.39879921e+04-5.57113251e+01-5.03717531e+00 8.30928098e-02-6.46761776e-05    3
 2.54418217e-08-3.97742990e-12-4.78544725e+04 5.00743814e+01                   4
MTBE-OO                 C   5H  11O   3     G    300.00   3500.00 1650.00      1
 1.64806414e+01 3.48147967e-02-1.47688703e-05 3.00165497e-09-2.41352085e-13    2
-3.59678543e+04-5.02874977e+01 2.84930338e+00 6.78604645e-02-4.48103865e-05    3
 1.51396413e-08-2.08044093e-12-3.14695128e+04 2.23020656e+01                   4
MTBE-QOOH               C   5H  11O   3     G    300.00   3500.00 1320.00      1
 1.54436168e+01 3.66620460e-02-1.53964709e-05 3.18866684e-09-2.64826231e-13    2
-2.86187066e+04-4.25445305e+01 1.39866731e+00 7.92224989e-02-6.37606219e-05    3
 2.76150057e-08-4.89102678e-12-2.49108399e+04 2.91135556e+01                   4
MTBE-OOQOOH             C   5H  11O   5     G    300.00   3500.00 1360.00      1
 1.70053290e+01 4.31260447e-02-1.99573142e-05 4.44658567e-09-3.89314825e-13    2
-4.64302953e+04-4.61328204e+01 4.65469144e+00 7.94514494e-02-6.00220987e-05    3
 2.40861860e-08-3.99953546e-12-4.30709219e+04 1.72494988e+01                   4
MTBE-OQOOH              C   5H  10O   4     G    300.00   3500.00 1750.00      1
 2.60727540e+01 2.16561806e-02-7.50837534e-06 1.18094342e-09-6.95948255e-14    2
-6.60762144e+04-1.03020563e+02 2.39248740e+00 7.57825044e-02-5.39023672e-05    3
 1.88548451e-08-2.59443792e-12-5.77881211e+04 2.44748864e+01                   4
MACRIL                  C   4H   6O   2     G    300.00   3500.00 1110.00      1
 9.14034170e+00 2.10870487e-02-7.42259201e-06 1.25044324e-09-8.33063961e-14    2
-4.12827790e+04-1.50267980e+01-1.13135759e+00 5.81021813e-02-5.74430415e-05    3
 3.12927552e-08-6.84959288e-12-3.90024617e+04 3.56001682e+01                   4
MCROT                   C   5H   8O   2     G    300.00   3500.00 1270.00      1
 1.13738844e+01 2.61318045e-02-8.74855270e-06 1.35831542e-09-8.00175424e-14    2
-4.63062145e+04-2.54801444e+01 2.72064698e-01 6.10981658e-02-5.00474046e-05    3
 2.30375028e-08-4.34757411e-12-4.34863523e+04 3.07332407e+01                   4
MB                      C   5H  10O   2     G    300.00   3500.00 1800.00      1
 1.24284215e+01 3.57133465e-02-1.61592897e-05 3.52094154e-09-3.02693558e-13    2
-6.07702345e+04-3.65220644e+01 2.77831323e+00 5.71580317e-02-3.40298606e-05    3
 1.01396715e-08-1.22196161e-12-5.72961955e+04 1.57063350e+01                   4
ALDEST                  C   6H  10O   3     G    300.00   3500.00 1800.00      1
 1.79608751e+01 3.27577411e-02-1.29904882e-05 2.50013886e-09-1.93431595e-13    2
-7.48983172e+04-5.99171164e+01 5.24137857e+00 6.10232889e-02-3.65451114e-05    3
 1.12240734e-08-1.40508916e-12-7.03192984e+04 8.92345209e+00                   4
UME7                    C   8H  14O   2     G    300.00   3500.00 1800.00      1
 2.58473881e+01 3.62113250e-02-1.33123979e-05 2.32937382e-09-1.61944423e-13    2
-5.91274202e+04-1.03960086e+02 2.21977770e+00 8.87171259e-02-5.70672320e-05    3
 1.85348679e-08-2.41270749e-12-5.06214805e+04 2.39174702e+01                   4
UME10                   C  11H  20O   2     G    300.00   3500.00 1800.00      1
 3.48566662e+01 5.08631766e-02-1.90027515e-05 3.39432409e-09-2.41664372e-13    2
-7.27334574e+04-1.48477352e+02 1.08700085e+00 1.25906877e-01-8.15391689e-05    3
 2.65559601e-08-3.45855827e-12-6.05763778e+04 3.42911218e+01                   4
MD                      C  11H  22O   2     G    300.00   3500.00 1800.00      1
 3.32942929e+01 6.02277988e-02-2.43433692e-05 4.77523343e-09-3.75629796e-13    2
-8.61538203e+04-1.40508544e+02 1.40263245e+00 1.31098155e-01-8.34019997e-05    3
 2.66488003e-08-3.41362519e-12-7.46728226e+04 3.20957753e+01                   4
C12H18                  C  12H  18          G    300.00   3500.00 1800.00      1
 8.44296021e+01 4.93170081e-02-2.86268137e-05 8.86979321e-09-1.00373559e-12    2
-8.94265355e+04-4.12065852e+02-1.18024932e+01 2.63166109e-01-2.06834398e-04    3
 7.48726021e-08-1.01707924e-11-5.47829811e+04 1.08762323e+02                   4
C12H22                  C  12H  22          G    300.00   3500.00 1760.00      1
 3.60687753e+01 4.93532020e-02-1.68932932e-05 2.64867330e-09-1.56935214e-13    2
-2.29291105e+04-1.58689916e+02-2.71855190e+00 1.37506218e-01-9.20237048e-05    3
 3.11071626e-08-4.19933426e-12-9.27597134e+03 5.03635283e+01                   4
ALDINS                  C  13H  20O   1     G    300.00   3500.00 1800.00      1
 8.44296021e+01 4.93170081e-02-2.86268137e-05 8.86979321e-09-1.00373559e-12    2
-8.94265355e+04-4.12065852e+02-1.18024932e+01 2.63166109e-01-2.06834398e-04    3
 7.48726021e-08-1.01707924e-11-5.47829811e+04 1.08762323e+02                   4
U2ME12                  C  13H  22O   2     G    300.00   3500.00 1610.00      1
 3.12799471e+01 7.15415825e-02-3.01181493e-05 6.08643057e-09-4.87334707e-13    2
-6.28268107e+04-1.24478604e+02 1.12650721e+00 1.46456961e-01-9.99150859e-05    3
 3.49878536e-08-4.97513331e-12-5.31174030e+04 3.53544123e+01                   4
UME16                   C  17H  32O   2     G    300.00   3500.00 1580.00      1
 4.52339567e+01 8.65152658e-02-3.05153568e-05 4.60675062e-09-2.26752937e-13    2
-9.22046801e+04-1.94026820e+02-6.34895688e+00 2.17104920e-01-1.54492877e-04    3
 5.69179405e-08-8.50383995e-12-7.59044794e+04 7.84262260e+01                   4
MPA                     C  17H  34O   2     G    300.00   3500.00 1570.00      1
 4.76347797e+01 8.91363204e-02-3.14080901e-05 4.73915928e-09-2.33379248e-13    2
-1.08404909e+05-2.13800468e+02-6.71212943e+00 2.27599783e-01-1.63698023e-04    3
 6.09132283e-08-9.17829469e-12-9.13399797e+04 7.29065183e+01                   4
MLIN1                   C  19H  32O   2     G    300.00   3500.00 1790.00      1
 6.02396150e+01 7.58945246e-02-2.57645421e-05 3.83449540e-09-2.03418694e-13    2
-7.74468643e+04-2.75096751e+02-2.53501003e+00 2.16173016e-01-1.43316351e-04    3
 4.76154297e-08-6.31807433e-12-5.49735486e+04 6.43028947e+01                   4
MLINO                   C  19H  34O   2     G    300.00   3500.00 1800.00      1
 6.05955634e+01 8.00185145e-02-2.72219283e-05 4.09058136e-09-2.22036704e-13    2
-9.16175349e+04-2.76065883e+02-1.22142713e+00 2.17389604e-01-1.41697837e-04    3
 4.64890659e-08-6.11071512e-12-6.93634183e+04 5.85005654e+01                   4
MEOLE                   C  19H  36O   2     G    300.00   3500.00 1800.00      1
 5.99430871e+01 8.58698870e-02-2.97676152e-05 4.64268484e-09-2.70021926e-13    2
-1.05323851e+05-2.71321302e+02-2.40329819e-02 2.19130154e-01-1.40817838e-04    3
 4.57723968e-08-5.98248192e-12-8.37356874e+04 5.32332617e+01                   4
MSTEA                   C  19H  38O   2     G    300.00   3500.00 1590.00      1
 5.57521905e+01 9.44092802e-02-3.21197954e-05 4.65296548e-09-2.12922090e-13    2
-1.17225838e+05-2.54579471e+02-7.52353585e+00 2.53593497e-01-1.82293585e-04    3
 6.76189151e-08-1.01132286e-11-9.71041567e+04 8.00324380e+01                   4
RMP3                    C   4H   7O   2     G    300.00   3500.00 1800.00      1
 9.46731366e+00 2.78903348e-02-1.31079832e-05 2.94998237e-09-2.60075468e-13    2
-3.18264559e+04-1.93081416e+01 3.67472849e+00 4.07627463e-02-2.38349927e-05    3
 6.92294888e-09-8.11876372e-13-2.97411253e+04 1.20425377e+01                   4
RMCROTA                 C   5H   7O   2     G    300.00   3500.00 1430.00      1
 1.57189270e+01 1.69463364e-02-4.46708471e-06 5.66631994e-10-2.76622249e-14    2
-3.23219578e+04-4.94508670e+01 1.47581648e-01 6.05025473e-02-5.01554178e-05    3
 2.18665542e-08-3.75142485e-12-2.78685530e+04 3.12413457e+01                   4
RMBX                    C   5H   9O   2     G    300.00   3500.00 1800.00      1
 1.54924675e+01 2.80794157e-02-1.20573290e-05 2.49322503e-09-2.04812831e-13    2
-3.97201853e+04-5.41810294e+01 2.13573336e+00 5.77610471e-02-3.67920218e-05    3
 1.16542224e-08-1.47717357e-12-3.49117610e+04 1.81084020e+01                   4
RALDEST                 C   6H   9O   3     G    300.00   3500.00 1800.00      1
 1.17688628e+01 4.16586301e-02-2.02330620e-05 4.68126733e-09-4.21941069e-13    2
-4.91007180e+04-2.27507760e+01 5.76645050e+00 5.49973242e-02-3.13486404e-05    3
 8.79814823e-09-9.93730082e-13-4.69398496e+04 9.73553178e+00                   4
RUME7                   C   8H  13O   2     G    300.00   3500.00 1800.00      1
 1.85903455e+01 4.63199612e-02-2.12076312e-05 4.67919509e-09-4.06994570e-13    2
-3.29183971e+04-6.07637962e+01 2.66158696e+00 8.17172025e-02-5.07053322e-05    3
 1.56042696e-08-1.92436602e-12-2.71840440e+04 2.54459681e+01                   4
RME7                    C   8H  15O   2     G    300.00   3500.00 1800.00      1
 2.40410389e+01 4.26053899e-02-1.71372003e-05 3.34440558e-09-2.61909736e-13    2
-4.89929734e+04-9.20931859e+01 2.93892074e+00 8.94989857e-02-5.62151968e-05    3
 1.78177376e-08-2.27209474e-12-4.13962109e+04 2.21158795e+01                   4
RUME10                  C  11H  19O   2     G    300.00   3500.00 1450.00      1
 2.35916391e+01 6.52041680e-02-2.68467493e-05 5.44034817e-09-4.42864583e-13    2
-3.58672712e+04-8.27430136e+01 1.64400787e+00 1.25749358e-01-8.94797041e-05    3
 3.42371090e-08-5.40782334e-12-2.95024582e+04 3.12965600e+01                   4
RMDX                    C  11H  21O   2     G    300.00   3500.00 1800.00      1
 2.51620787e+01 7.14154782e-02-3.28251105e-05 7.27502335e-09-6.35223044e-13    2
-5.95987228e+04-9.23572152e+01 1.85440069e+00 1.23210318e-01-7.59874772e-05    3
 2.32610851e-08-2.85550940e-12-5.12079587e+04 3.37888005e+01                   4
RUME16                  C  17H  31O   2     G    300.00   3500.00 1790.00      1
 5.62816136e+01 7.14355326e-02-2.43271963e-05 3.65698891e-09-1.98260059e-13    2
-7.53410003e+04-2.53924454e+02 9.94523443e-01 1.94982103e-01-1.27857842e-04    3
 4.22158885e-08-5.58358123e-12-5.55482221e+04 4.49928047e+01                   4
RMPAX                   C  17H  33O   2     G    300.00   3500.00 1570.00      1
 4.65991995e+01 8.79958434e-02-3.11818055e-05 4.72866732e-09-2.34133595e-13    2
-8.86750545e+04-2.03460515e+02-5.53001449e+00 2.20809128e-01-1.58073478e-04    3
 5.86104816e-08-8.81404033e-12-7.23064813e+04 7.15470262e+01                   4
RMLIN1X                 C  19H  31O   2     G    300.00   3500.00 1800.00      1
 5.95150805e+01 7.42460884e-02-2.53824685e-05 3.82833284e-09-2.08614183e-13    2
-4.82863792e+04-2.69048888e+02-9.12525139e-01 2.08529657e-01-1.37285442e-04    3
 4.52738785e-08-5.96493998e-12-2.65324412e+04 5.79979195e+01                   4
RMLIN1A                 C  19H  31O   2     G    300.00   3500.00 1800.00      1
 5.95150805e+01 7.42460884e-02-2.53824685e-05 3.82833284e-09-2.08614183e-13    2
-4.82863792e+04-2.69048888e+02-9.12525139e-01 2.08529657e-01-1.37285442e-04    3
 4.52738785e-08-5.96493998e-12-2.65324412e+04 5.79979195e+01                   4
RMLINA                  C  19H  33O   2     G    300.00   3500.00 1800.00      1
 5.71954572e+01 8.40022526e-02-3.15645609e-05 5.64020282e-09-4.00097416e-13    2
-6.69574792e+04-2.54485524e+02-1.30856007e+00 2.14011180e-01-1.39905334e-04    3
 4.57664149e-08-5.97318243e-12-4.58960330e+04 6.21504214e+01                   4
RMLINX                  C  19H  33O   2     G    300.00   3500.00 1800.00      1
 5.71954572e+01 8.40022526e-02-3.15645609e-05 5.64020282e-09-4.00097416e-13    2
-6.69574792e+04-2.54485524e+02-1.30856007e+00 2.14011180e-01-1.39905334e-04    3
 4.57664149e-08-5.97318243e-12-4.58960330e+04 6.21504214e+01                   4
RMEOLES                 C  19H  35O   2     G    300.00   3500.00 1800.00      1
 5.65771897e+01 8.98806670e-02-3.42288637e-05 6.24737169e-09-4.55217496e-13    2
-8.06885314e+04-2.49965187e+02-1.57103417e-01 2.15956874e-01-1.39292369e-04    3
 4.51597812e-08-5.85971882e-12-6.02641859e+04 5.70926426e+01                   4
RMEOLEA                 C  19H  35O   2     G    300.00   3500.00 1800.00      1
 5.65771897e+01 8.98806670e-02-3.42288637e-05 6.24737169e-09-4.55217496e-13    2
-8.06885314e+04-2.49965187e+02-1.57103417e-01 2.15956874e-01-1.39292369e-04    3
 4.51597812e-08-5.85971882e-12-6.02641859e+04 5.70926426e+01                   4
RSTEAX                  C  19H  37O   2     G    300.00   3500.00 1590.00      1
 5.46335770e+01 9.34230794e-02-3.19964368e-05 4.67181990e-09-2.16707128e-13    2
-9.74617250e+04-2.43777070e+02-6.34709276e+00 2.46833569e-01-1.76723314e-04    3
 6.53539487e-08-9.75792235e-12-7.80698720e+04 7.86982222e+01                   4
ETMB583                 C   5H   8O   3     G    300.00   3500.00 1270.00      1
 1.75630364e+01 2.35383861e-02-7.56913212e-06 1.05837473e-09-4.95698456e-14    2
-6.27369638e+04-6.15054251e+01-4.60165687e+00 9.33484435e-02-9.00219558e-05    3
 4.43406969e-08-8.56971200e-12-5.71071317e+04 5.07241436e+01                   4
KEHYMB                  C   5H   8O   5     G    300.00   3500.00 1200.00      1
 1.28585854e+01 3.05267696e-02-1.05263783e-05 1.70287730e-09-1.06411275e-13    2
-6.04915273e+04-3.42459470e+01-2.28352155e+00 8.10004595e-02-7.36184906e-05    3
 3.67540508e-08-7.40873909e-12-5.68574216e+04 4.15666987e+01                   4
C7H15COCHO              C   9H  16O   2     G    300.00   3500.00 1780.00      1
 3.02051070e+01 3.84107404e-02-1.30453988e-05 2.02881282e-09-1.19347924e-13    2
-6.67956482e+04-1.25747099e+02 3.59041212e-01 1.05480551e-01-6.95649021e-05    3
 2.31971661e-08-3.09243126e-12-5.61704488e+04 3.54525564e+01                   4
ALD9                    C   9H  18O   1     G    300.00   3500.00 1140.00      1
 1.64741951e+01 5.58925365e-02-1.69806972e-05 1.83483646e-09-1.30758059e-14    2
-4.58697504e+04-4.72673092e+01-2.96684223e+00 1.24106702e-01-1.06736179e-04    3
 5.43234221e-08-1.15237306e-11-4.14371939e+04 4.90717830e+01                   4
MEALD9                  C  10H  18O   3     G    300.00   3500.00  990.00      1
 2.52719799e+01 4.25885173e-02 2.29436427e-06-6.10865001e-09 1.00091979e-12    2
-8.74828172e+04-8.25654359e+01-5.97961626e+00 1.68857593e-01-1.89022416e-04    3
 1.22724199e-07-3.15326279e-11-8.12950012e+04 6.78913613e+01                   4
ETEROMD                 C  11H  20O   3     G    300.00   3500.00 1760.00      1
 4.14249232e+01 4.51122010e-02-1.56530058e-05 2.49213985e-09-1.50324644e-13    2
-8.95581286e+04-1.84296556e+02-1.24328084e-01 1.39542318e-01-9.61332188e-05    3
 3.29770690e-08-4.48057027e-12-7.49327921e+04 3.96429290e+01                   4
MDKETO                  C  11H  20O   5     G    300.00   3500.00 1420.00      1
 2.98411849e+01 7.16595757e-02-3.12595602e-05 6.71204679e-09-5.73522213e-13    2
-1.08207341e+05-1.07784029e+02 3.72296288e+00 1.45232032e-01-1.08976944e-04    3
 4.31990813e-08-6.99729589e-12-1.00789766e+05 2.73798286e+01                   4
MEALDU12                C  13H  22O   3     G    300.00   3500.00 1070.00      1
 2.71187290e+01 6.80017640e-02-1.53844386e-05-3.62279043e-10 3.31896805e-13    2
-8.26297086e+04-8.79500630e+01-7.00276451e+00 1.95558749e-01-1.94202642e-04    3
 1.11050932e-07-2.56992272e-11-7.53277090e+04 7.89750333e+01                   4
ETEROMPA                C  17H  32O   3     G    300.00   3500.00 1310.00      1
 4.32126688e+01 9.17256515e-02-3.02788110e-05 4.53882530e-09-2.50045062e-13    2
-1.06117741e+05-1.75617614e+02-8.73011642e+00 2.50329576e-01-2.11886358e-04    3
 9.69599687e-08-1.78876679e-11-9.25087311e+04 8.90022604e+01                   4
KHMLIN1                 C  19H  30O   5     G    300.00   3500.00 1690.00      1
 6.18941876e+01 8.22994971e-02-3.10180831e-05 5.38913501e-09-3.62607369e-13    2
-9.79974619e+04-2.72277440e+02-3.09268632e+00 2.36114583e-01-1.67540349e-04    3
 5.92440722e-08-8.32931406e-12-7.60318985e+04 7.53471279e+01                   4
MLIN1OOH                C  19H  34O   4     G    300.00   3500.00 1800.00      1
 6.05955634e+01 8.00185145e-02-2.72219283e-05 4.09058136e-09-2.22036704e-13    2
-9.16175349e+04-2.76065883e+02-1.22142713e+00 2.17389604e-01-1.41697837e-04    3
 4.64890659e-08-6.11071512e-12-6.93634183e+04 5.85005654e+01                   4
MLINOOH                 C  19H  36O   4     G    300.00   3500.00 1800.00      1
 6.05955634e+01 8.00185145e-02-2.72219283e-05 4.09058136e-09-2.22036704e-13    2
-9.16175349e+04-2.76065883e+02-1.22142713e+00 2.17389604e-01-1.41697837e-04    3
 4.64890659e-08-6.11071512e-12-6.93634183e+04 5.85005654e+01                   4
MSTEAKETO               C  19H  36O   5     G    300.00   3500.00 1630.00      1
 6.13348278e+01 9.80436835e-02-3.77033626e-05 6.80816985e-09-4.83388138e-13    2
-1.42870187e+05-2.70834379e+02-4.17722885e-01 2.49583685e-01-1.77157352e-04    3
 6.38445663e-08-9.23130171e-12-1.22738855e+05 5.72570440e+01                   4
RMBOOX                  C   5H   9O   4     G    300.00   3500.00 1350.00      1
 2.46557077e+01 1.60203217e-02-2.33017820e-06-2.09433435e-10 5.96257322e-14    2
-5.87318869e+04-9.28197899e+01-3.02577563e+00 9.80395314e-02-9.34626335e-05    3
 4.47942482e-08-8.27438938e-12-5.12578864e+04 4.90347058e+01                   4
QMBOOX                  C   5H   9O   4     G    300.00   3500.00 1350.00      1
 2.46557077e+01 1.60203217e-02-2.33017820e-06-2.09433435e-10 5.96257322e-14    2
-5.87318869e+04-9.28197899e+01-3.02577563e+00 9.80395314e-02-9.34626335e-05    3
 4.47942482e-08-8.27438938e-12-5.12578864e+04 4.90347058e+01                   4
ZMBOOX                  C   5H   9O   6     G    300.00   3500.00 1310.00      1
 2.94016989e+01 1.57346327e-02-2.10564640e-06-2.30313524e-10 5.80532439e-14    2
-7.03637127e+04-1.09596866e+02-1.66570926e+00 1.10596948e-01-1.10726618e-04    3
 5.50475345e-08-1.04911544e-11-6.22240518e+04 4.86744631e+01                   4
QMDOOH                  C  11H  21O   4     G    300.00   3500.00 1800.00      1
 3.77681893e+01 6.05584615e-02-2.66377187e-05 5.63138780e-09-4.71383164e-13    2
-7.68263337e+04-1.55143434e+02 4.12866787e+00 1.35312954e-01-8.89331288e-05    3
 2.87037619e-08-3.67587957e-12-6.47161059e+04 2.69206740e+01                   4
RMDOOX                  C  11H  21O   4     G    300.00   3500.00 1800.00      1
 3.96894066e+01 5.38224995e-02-2.02774959e-05 3.64793757e-09-2.61216218e-13    2
-8.38472353e+04-1.67546754e+02 4.70466734e+00 1.31566364e-01-8.50640501e-05    3
 2.76429576e-08-3.59385789e-12-7.12527292e+04 2.17979534e+01                   4
ZMDOOH                  C  11H  21O   6     G    300.00   3500.00 1780.00      1
 4.89601112e+01 4.69646638e-02-1.61477787e-05 2.58757397e-09-1.58080064e-13    2
-9.96313670e+04-2.11226525e+02 6.91495065e+00 1.41448171e-01-9.57687114e-05    3
 3.24081480e-08-4.34636293e-12-8.46632899e+04 1.58608718e+01                   4
QMPAOOH                 C  17H  33O   4     G    300.00   3500.00 1800.00      1
 3.77681893e+01 6.05584615e-02-2.66377187e-05 5.63138780e-09-4.71383164e-13    2
-7.68263337e+04-1.55143434e+02 4.12866787e+00 1.35312954e-01-8.89331288e-05    3
 2.87037619e-08-3.67587957e-12-6.47161059e+04 2.69206740e+01                   4
RMPAOOX                 C  17H  33O   4     G    300.00   3500.00 1800.00      1
 3.96894066e+01 5.38224995e-02-2.02774959e-05 3.64793757e-09-2.61216218e-13    2
-8.38472353e+04-1.67546754e+02 4.70466734e+00 1.31566364e-01-8.50640501e-05    3
 2.76429576e-08-3.59385789e-12-7.12527292e+04 2.17979534e+01                   4
ZMPAOOH                 C  17H  33O   6     G    300.00   3500.00 1780.00      1
 4.89601112e+01 4.69646638e-02-1.61477787e-05 2.58757397e-09-1.58080064e-13    2
-9.96313670e+04-2.11226525e+02 6.91495065e+00 1.41448171e-01-9.57687114e-05    3
 3.24081480e-08-4.34636293e-12-8.46632899e+04 1.58608718e+01                   4
HEXENAL                 C   6H  10O   1     G    300.00   3500.00 1800.00      1
 2.52910440e+01 1.04447230e-02 8.54445711e-07-1.11418266e-09 1.52698388e-13    2
-2.77614674e+04-1.05594851e+02-9.42771449e-01 6.87420906e-02-4.77266940e-05    3
 1.68788320e-08-2.34633143e-12-1.83172939e+04 3.63880312e+01                   4
QMLIN1OOX               C  19H  31O   4     G    300.00   3500.00 1610.00      1
 5.66825592e+01 9.03049049e-02-3.59434729e-05 6.72610645e-09-4.95506472e-13    2
-6.74923705e+04-2.44601807e+02-2.71828944e+00 2.37884653e-01-1.73440133e-04    3
 6.36605411e-08-9.33625720e-12-4.83652972e+04 7.02616646e+01                   4
RMLIN1OOX               C  19H  31O   4     G    300.00   3500.00 1650.00      1
 5.48798838e+01 9.05843890e-02-3.54321228e-05 6.50176129e-09-4.69049126e-13    2
-7.13229385e+04-2.34809026e+02-1.47497533e+00 2.27202229e-01-1.59630160e-04    3
 5.66827862e-08-8.07223473e-12-5.27258349e+04 6.52917144e+01                   4
ZMLIN1OOX               C  19H  31O   6     G    300.00   3500.00 1690.00      1
 6.61919906e+01 8.18444488e-02-3.03706310e-05 5.17171901e-09-3.39001412e-13    2
-8.83104234e+04-2.93138165e+02 7.95448659e-01 2.36629163e-01-1.67753514e-04    3
 5.93661501e-08-8.35592908e-12-6.62063922e+04 5.66777785e+01                   4
RMLIN1OH                C  19H  33O   3     G    300.00   3500.00 1800.00      1
 8.28450490e+01 6.90025877e-02-5.05706431e-05 1.59456839e-08-1.77055095e-12    2
-1.00000197e+05-4.01748327e+02-1.67494614e+01 2.90323722e-01-2.35004922e-04    3
 8.42546759e-08-1.12579110e-11-6.41461731e+04 1.37277939e+02                   4
QMLINOOX                C  19H  33O   4     G    300.00   3500.00 1760.00      1
 6.81310039e+01 7.45379717e-02-2.47877879e-05 3.55693193e-09-1.75306750e-13    2
-8.29474487e+04-3.08878588e+02 1.76450133e-02 2.29341060e-01-1.56722238e-04    3
 5.35321025e-08-7.27405257e-12-5.89715464e+04 5.82344177e+01                   4
RMLINOOX                C  19H  33O   4     G    300.00   3500.00 1780.00      1
 6.32132488e+01 8.05239268e-02-2.78197685e-05 4.27200551e-09-2.39927626e-13    2
-8.77238934e+04-2.82700435e+02 1.99661291e+00 2.18089401e-01-1.43745730e-04    3
 4.76899685e-08-6.33795613e-12-6.59307710e+04 4.79327766e+01                   4
RMLIN1OHOO              C  19H  33O   5     G    300.00   3500.00 1120.00      1
 4.66382276e+01 9.44918900e-02-2.04259617e-05-5.03856990e-10 4.25993739e-13    2
-9.66680676e+04-1.74384019e+02-1.26774253e+01 3.06333507e-01-3.04142414e-04    3
 1.68374983e-07-3.72701760e-11-8.33813614e+04 1.18501883e+02                   4
ZMLINOOX                C  19H  33O   6     G    300.00   3500.00 1530.00      1
 6.14087103e+01 8.58331760e-02-2.98017545e-05 4.63939550e-09-2.65660848e-13    2
-9.65914219e+04-2.81173972e+02 1.31186641e+00 2.42949108e-01-1.83836982e-04    3
 7.17571416e-08-1.12326128e-11-7.82017876e+04 3.43158093e+01                   4
RMEOLEOOX               C  19H  35O   4     G    300.00   3500.00 1800.00      1
 5.68288338e+01 9.87024759e-02-3.87236377e-05 7.19531818e-09-5.31280167e-13    2
-1.23280982e+05-2.44956703e+02 2.29714005e+00 2.19884018e-01-1.39708256e-04    3
 4.45970286e-08-5.72596217e-12-1.03649572e+05 5.01801999e+01                   4
QMEOLEOOH               C  19H  35O   4     G    300.00   3500.00 1800.00      1
 6.66288155e+01 8.44466821e-02-2.89700531e-05 4.40901581e-09-2.44933389e-13    2
-1.50877975e+05-3.00441870e+02-9.98788075e-01 2.34730246e-01-1.54206356e-04    3
 5.07928317e-08-6.68713004e-12-1.26532038e+05 6.55728279e+01                   4
ZMEOLEOOX               C  19H  35O   6     G    300.00   3500.00 1540.00      1
 5.74950069e+01 9.92606520e-02-3.35004160e-05 5.08063928e-09-2.82240577e-13    2
-1.09648464e+05-2.38315332e+02 2.38451835e+00 2.42404778e-01-1.72926513e-04    3
 6.54382570e-08-1.00805551e-11-9.26744334e+04 5.13566581e+01                   4
RMEOLEOH                C  19H  37O   3     G    300.00   3500.00 1800.00      1
 8.79849800e+01 7.07215853e-02-4.99029476e-05 1.57162432e-08-1.74835864e-12    2
-1.30787157e+05-4.30015035e+02-1.57729922e+01 3.01294857e-01-2.42047341e-04    3
 8.68808331e-08-1.16323295e-11-9.34342873e+04 1.31544755e+02                   4
QMSTEAOOH               C  19H  37O   4     G    300.00   3500.00 1230.00      1
-1.30612119e+02 6.00365428e-01-4.85197524e-04 1.58690699e-07-1.80918285e-11    2
 1.24045733e+04 7.12083772e+02 2.15554530e+01 1.05511534e-01 1.18282834e-04    3
-1.68398926e-07 4.83898026e-11-2.50286495e+04-5.35376471e+01                   4
RMSTEAOOX               C  19H  37O   4     G    300.00   3500.00 1250.00      1
-1.20700823e+02 5.67736642e-01-4.52750601e-04 1.47317718e-07-1.67528749e-11    2
 1.02039723e+04 6.60023999e+02 1.91170962e+01 1.20319300e-01 8.41502093e-05    3
-1.39029381e-07 4.05165449e-11-2.47505076e+04-4.57161070e+01                   4
RMEOLEOHOO              C  19H  37O   5     G    300.00   3500.00 1070.00      1
 4.98703764e+01 9.32941337e-02-1.10712954e-05-4.86534745e-09 9.98405301e-13    2
-1.26041658e+05-1.89643846e+02-1.31696044e+01 3.28957613e-01-3.41440659e-04    3
 2.00972262e-07-4.70944942e-11-1.12551102e+05 1.18752821e+02                   4
ZMSTEAOOH               C  19H  37O   6     G    300.00   3500.00 1250.00      1
-6.22995272e+01 3.41575939e-01-2.69706989e-04 8.71969158e-08-9.87435428e-12    2
 1.57160046e+04 3.57020389e+02 1.61954270e+01 9.03920855e-02 3.17136355e-05    3
-7.35607505e-08 2.22771790e-11-3.90773394e+03-3.91880335e+01                   4
NO                      N   1O   1          G    200.00   3500.00  800.00      1
 2.84621514e+00 2.06354049e-03-1.06904718e-06 2.65706534e-10-2.54948690e-14    2
 1.00671113e+04 8.61842850e+00 4.25026595e+00-4.95671355e-03 1.20939291e-05    3
-1.07034404e-08 3.40236355e-12 9.84246312e+03 2.15799985e+00                   4
N2O                     N   2O   1          G    200.00   3500.00 1420.00      1
 4.85543737e+00 2.58052405e-03-9.33593927e-07 1.54088379e-10-9.24861941e-15    2
 8.05595822e+03-2.39060931e+00 2.51620680e+00 9.16990594e-03-7.89420860e-06    3
 3.42198259e-09-5.84582107e-13 8.72029970e+03 9.71509326e+00                   4
NO2                     N   1O   2          G    200.00   3500.00 1800.00      1
 4.19813812e+00 3.78881343e-03-2.08225979e-06 5.53837903e-10-5.45690310e-14    2
 2.49824361e+03 3.49647478e+00 2.86592220e+00 6.74929324e-03-4.54932631e-06    3
 1.46756624e-09-1.81475745e-13 2.97784134e+03 1.07067052e+01                   4
HNO                     H   1N   1O   1     G    200.00   3500.00  700.00      1
 2.88552847e+00 3.71507602e-03-9.89194593e-07 1.60505686e-10-1.61198707e-14    2
 1.18465422e+04 9.10108579e+00 4.47186924e+00-5.34972841e-03 1.84353863e-05    3
-1.83390952e-08 6.59088044e-12 1.16244545e+04 2.01371655e+00                   4
HNO2                    H   1N   1O   2     G    200.00   3500.00  700.00      1
 1.72007297e+00 1.13464166e-02-6.67663346e-06 1.82835452e-09-1.88889112e-13    2
-6.26025905e+03 1.58192354e+01 3.09881790e+00 3.46787417e-03 1.02059575e-05    3
-1.42503035e-08 5.55348876e-12-6.45328334e+03 9.65935184e+00                   4
HONO                    H   1N   1O   2     G    200.00   3500.00 1450.00      1
 5.99816573e+00 3.29505590e-03-1.07588917e-06 1.49768801e-10-6.76019245e-15    2
-1.16909496e+04-5.24156231e+00 2.71684795e+00 1.23469670e-02-1.04399352e-05    3
 4.45507730e-09-7.49054762e-13-1.07393674e+04 1.18081173e+01                   4
HONO2                   H   1N   1O   3     G    200.00   3500.00 1480.00      1
 8.72243727e+00 3.29016335e-03-9.97287988e-07 9.83681568e-11 7.21043264e-16    2
-1.96262632e+04-2.01737933e+01 1.12599201e+00 2.38210965e-02-2.18056662e-05    3
 9.47151148e-09-1.58258019e-12-1.73777154e+04 1.94527902e+01                   4
N2H2                    N   2H   2          G    200.00   3500.00  700.00      1
 1.61507707e+00 8.37729344e-03-2.70267456e-06 3.47805161e-10-1.28897270e-14    2
 2.32788099e+04 1.47543853e+01 4.76517120e+00-9.62324442e-03 3.58699066e-05    3
-3.63879864e-08 1.31070358e-11 2.28377967e+04 6.80561701e-01                   4
H2NN                    N   2H   2          G    200.00   3500.00  700.00      1
 1.58440836e+00 9.29486031e-03-4.50990678e-06 1.06229464e-09-9.86121908e-14    2
 3.53712259e+04 1.46993890e+01 4.53650989e+00-7.57429125e-03 3.16382751e-05    3
-3.33645453e-08 1.21966878e-11 3.49579317e+04 1.51014624e+00                   4
HNNO                    H   1O   1N   2     G    300.00   3500.00 1360.00      1
 4.88500313e+00 5.60936882e-03-2.60717813e-06 5.93838981e-10-5.41495052e-14    2
 2.58926738e+04 6.01979772e-01 2.29344827e+00 1.32315890e-02-1.10140386e-05    3
 4.71484903e-09-8.11688117e-13 2.65975767e+04 1.39015974e+01                   4
NH2NO                   N   2H   2O   1     G    300.00   3500.00 1800.00      1
 5.77099677e+00 9.34065649e-03-4.91078058e-06 1.15317940e-09-1.04142547e-13    2
 6.27743926e+03-6.42401937e+00 1.47077488e+00 1.88967051e-02-1.28741545e-05    3
 4.10257713e-09-5.13781121e-13 7.82551914e+03 1.68496786e+01                   4
NH2OH                   N   1H   3O   1     G    200.00   3500.00 1140.00      1
 3.89950467e+00 8.10759734e-03-2.78780456e-06 4.26313819e-10-2.40531623e-14    2
-6.86348420e+03 3.69890799e+00 2.36719772e+00 1.34841130e-02-9.86216723e-06    3
 4.56336801e-09-9.31301888e-13-6.51411822e+03 1.12921788e+01                   4
HNOH                    H   2N   1O   1     G    200.00   3500.00 1800.00      1
 3.80328695e+00 5.45108884e-03-2.14629755e-06 4.23543084e-10-3.43983592e-14    2
 1.05861530e+04 4.48881970e+00 2.57438368e+00 8.18198500e-03-4.42204435e-06    3
 1.26641227e-09-1.51463524e-13 1.10285582e+04 1.11399006e+01                   4
NH3                     H   3N   1          G    200.00   3500.00  700.00      1
 2.51781806e+00 5.95384020e-03-2.00551772e-06 3.21049849e-10-1.88806092e-14    2
-6.46278678e+03 7.18902507e+00 4.05091143e+00-2.80669335e-03 1.67670542e-05    3
-1.75575900e-08 6.36634792e-12-6.67741985e+03 3.39551759e-01                   4
N2H4                    N   2H   4          G    200.00   3500.00 1780.00      1
 6.33303400e+00 6.50860326e-03-1.68647151e-06 1.37723180e-10 3.10853742e-15    2
 8.61374390e+03-1.06617456e+01 1.71754273e+00 1.68804937e-02-1.04268287e-05    3
 3.41126518e-09-4.56658598e-13 1.02568588e+04 1.42666857e+01                   4
N                       N   1               G    200.00   3500.00 1800.00      1
 2.42215558e+00 1.52655400e-04-9.87414140e-08 2.32518157e-11-1.22034408e-15    2
 5.61344053e+04 4.62162565e+00 2.50554288e+00-3.26497066e-05 5.56795078e-08    3
-3.39411183e-11 6.72311898e-15 5.61043859e+04 4.17031620e+00                   4
NO3                     N   1O   3          G    200.00   3500.00 1380.00      1
 7.84336716e+00 1.94266710e-03-6.08796317e-07 6.42441728e-11-1.29683643e-16    2
 5.97435401e+03-1.61838239e+01 7.80027972e-01 2.24161140e-02-2.28625430e-05    3
 1.08148464e-08-1.94770256e-12 7.92383562e+03 2.01676897e+01                   4
NH                      N   1H   1          G    200.00   3500.00 1670.00      1
 2.48662851e+00 1.81565419e-03-7.12540990e-07 1.51936822e-10-1.23899396e-14    2
 4.24864648e+04 7.43461481e+00 3.66298285e+00-1.00196100e-03 1.81825110e-06    3
-8.58359421e-10 1.38852013e-13 4.20935624e+04 1.15612280e+00                   4
NNH                     N   2H   1          G    200.00   3500.00  740.00      1
 2.70691636e+00 4.73245705e-03-2.26389308e-06 5.23129607e-10-4.76635083e-14    2
 2.90245413e+04 1.03117271e+01 4.29167557e+00-3.83380896e-03 1.51001596e-05    3
-1.51201611e-08 5.23723201e-12 2.87899969e+04 3.14335908e+00                   4
NH2                     N   1H   2          G    200.00   3500.00 1280.00      1
 2.55273405e+00 3.54675616e-03-1.12718101e-06 1.61534558e-10-6.97198096e-15    2
 2.15912602e+04 8.13032049e+00 4.10678626e+00-1.30965699e-03 4.56392815e-06    3
-2.80258479e-09 5.71957580e-13 2.11934228e+04 2.49283473e-01                   4
H2NO                    N   1H   2O   1     G    200.00   3500.00  700.00      1
 2.72801503e+00 7.40936634e-03-3.46220932e-06 8.08344176e-10-7.54853132e-14    2
 6.86495538e+03 9.84388857e+00 3.66110547e+00 2.07742096e-03 7.96338790e-06    3
-1.00731770e-08 3.81077225e-12 6.73432272e+03 5.67507655e+00                   4
N2H3                    N   2H   3          G    200.00   3500.00 1800.00      1
 4.54460731e+00 6.62772188e-03-2.15038331e-06 3.20318484e-10-1.81983596e-14    2
 2.50493361e+04-4.68131456e-02 2.12003672e+00 1.20156565e-02-6.64032885e-06    3
 1.98326127e-09-2.49162636e-13 2.59221815e+04 1.30754687e+01                   4
HCN                     H   1C   1N   1     G    200.00   3500.00  780.00      1
 3.49786303e+00 3.76915263e-03-1.51027198e-06 3.01080795e-10-2.43629344e-14    2
 1.43955802e+04 3.23683725e+00 2.24572678e+00 1.01903642e-02-1.38587557e-05    3
 1.08553404e-08-3.40713845e-12 1.45909135e+04 8.96656338e+00                   4
HNC                     H   1N   1C   1     G    200.00   3500.00  700.00      1
 4.41179648e+00 2.12707772e-03-4.71967938e-07 1.02350842e-12 7.69770549e-15    2
 2.16589079e+04-1.07356900e+00 2.73172549e+00 1.17274834e-02-2.10442658e-05    3
 1.95936882e-08-6.98968253e-12 2.18941178e+04 6.43256315e+00                   4
HNCO                    H   1N   1C   1O   1G    200.00   3500.00 1050.00      1
 4.68274050e+00 5.27517072e-03-2.30255431e-06 4.91740878e-10-4.20405782e-14    2
-1.59709573e+04 2.61732213e-01 2.23902626e+00 1.45845583e-02-1.56016795e-05    3
 8.93562986e-09-2.05249034e-12-1.54577773e+04 1.21704701e+01                   4
HCNO                    H   1N   1C   1O   1G    200.00   3500.00  780.00      1
 4.79767989e+00 6.41431464e-03-3.21741500e-06 7.84733950e-10-7.49876248e-14    2
 1.84217969e+04-2.20789655e+00 6.69823249e-01 2.75828103e-02-4.39260604e-05    3
 3.55784480e-08-1.12268190e-11 1.90657425e+04 1.66810128e+01                   4
HOCN                    H   1N   1C   1O   1G    200.00   3500.00 1260.00      1
 5.08605511e+00 4.40745631e-03-1.67135012e-06 3.00184368e-10-2.12769812e-14    2
-3.69516510e+03-1.53122302e+00 2.95277826e+00 1.11797637e-02-9.73362087e-06    3
 4.56593609e-09-8.67656291e-13-3.15757934e+03 9.25362986e+00                   4
CH2NO                   C   1H   2N   1O   1G    200.00   3500.00 1800.00      1
 3.20402861e+00-6.01465229e-03 5.38459555e-05-6.82208900e-08 2.71923019e-11    2
 2.61694731e+04 1.15885287e+01 8.41613768e+00-1.75971169e-02 6.34980094e-05    3
-7.17957248e-08 2.76888067e-11 2.42931138e+04-1.66204929e+01                   4
CH3NO                   C   1H   3N   1O   1G    200.00   3500.00  700.00      1
 1.71612023e+00 1.65151446e-02-8.81735213e-06 2.26713782e-09-2.25490386e-13    2
 7.35980363e+03 1.71612002e+01 4.07025668e+00 3.06293627e-03 2.00088085e-05    3
-2.51863485e-08 9.57932617e-12 7.03022453e+03 6.64351414e+00                   4
CH3NO2                  C   1H   3N   1O   2G    200.00   3500.00 1800.00      1
 5.69934702e+00 1.38065590e-02-6.43453198e-06 1.45264650e-09-1.30225174e-13    2
-1.27635734e+04-5.01015454e+00 5.58676745e-01 2.52302708e-02-1.59542918e-05    3
 4.97848345e-09-6.19924750e-13-1.09129321e+04 2.28122254e+01                   4
CH3ONO                  C   1H   3O   2N   1G    200.00   3500.00  700.00      1
 2.81666880e+00 1.89749543e-02-1.04049678e-05 2.71704311e-09-2.72624825e-13    2
-9.44747973e+03 1.52094758e+01 5.07409813e+00 6.07535809e-03 1.72370239e-05    3
-2.36086633e-08 9.12941320e-12-9.76351983e+03 5.12385272e+00                   4
CH3ONO2                 C   1H   3N   1O   3G    200.00   3500.00 1800.00      1
 1.20582349e+01 7.66565964e-03-2.49975720e-06 3.22040139e-10-1.19528323e-14    2
-2.00738855e+04-3.71551232e+01 2.05585065e+00 2.98931803e-02-2.10226911e-05    3
 7.18238602e-09-9.64778650e-13-1.64730272e+04 1.69798673e+01                   4
CH3CN                   C   2H   3N   1     G    200.00   3500.00  700.00      1
 2.04918661e+00 1.63166629e-02-8.45703412e-06 2.11771923e-09-2.06450504e-13    2
 7.64801687e+03 1.30927477e+01 3.05185732e+00 1.05871160e-02 3.82056642e-06    3
-9.57523366e-09 3.96960410e-12 7.50764297e+03 8.61306859e+00                   4
CN                      C   1N   1          G    200.00   3500.00  890.00      1
 2.80498941e+00 1.99013252e-03-1.04863797e-06 2.95566175e-10-3.14165351e-14    2
 5.18669927e+04 7.89927659e+00 3.76469137e+00-2.32313471e-03 6.22091354e-06    3
-5.14979077e-09 1.49817811e-12 5.16961658e+04 3.38110713e+00                   4
NCN                     C   1N   2          G    200.00   3500.00 1540.00      1
 6.26178526e+00 8.14604797e-04-6.32168539e-08-5.68978404e-11 1.02757847e-14    2
 5.13388448e+04-9.55046093e+00 2.82367216e+00 9.74476868e-03-8.76142843e-06    3
 3.70856172e-09-6.01000118e-13 5.23977836e+04 8.52096413e+00                   4
NCO                     N   1C   1O   1     G    200.00   3500.00 1630.00      1
 5.49723477e+00 1.70371882e-03-5.14810248e-07 5.30241383e-11-1.05681650e-16    2
 1.33777864e+04-4.53940107e+00 2.90100728e+00 8.07482924e-03-6.37779530e-06    3
 2.45097304e-09-3.67889255e-13 1.42241566e+04 9.25436072e+00                   4
HNCN                    C   1H   1N   2     G    200.00   3500.00 1460.00      1
 5.71563451e+00 3.59039495e-03-1.19666866e-06 1.72409879e-10-8.44529375e-15    2
 3.58827350e+04-4.39973242e+00 3.04255634e+00 1.09138968e-02-8.72081438e-06    3
 3.60809286e-09-5.96747173e-13 3.66632738e+04 9.50791473e+00                   4
H2CN                    C   1H   2N   1     G    200.00   3500.00  700.00      1
 2.09516104e+00 9.19258717e-03-4.75958103e-06 1.19375089e-09-1.16674695e-13    2
 2.77113212e+04 1.25272169e+01 3.31830756e+00 2.20317847e-03 1.02177233e-05    3
-1.30703485e-08 4.97764652e-12 2.75400807e+04 7.06250770e+00                   4
HCNH                    C   1H   2N   1     G    200.00   3500.00  700.00      1
 2.20517224e+00 9.23158578e-03-4.92876098e-06 1.27407702e-09-1.27539972e-13    2
 3.17668288e+04 1.24496856e+01 2.93126391e+00 5.08249052e-03 3.96215742e-06    3
-7.19346431e-09 2.89658193e-12 3.16651760e+04 9.20569168e+00                   4
C2N2                    C   2N   2          G    200.00   3500.00  700.00      1
 5.66789418e+00 5.81681884e-03-2.89262860e-06 6.98368893e-10-6.54524579e-14    2
 3.52445641e+04-4.84945646e+00 2.74684240e+00 2.25085433e-02-3.86606096e-05    3
 3.47631127e-08-1.22314324e-11 3.56535113e+04 8.20106387e+00                   4
CH2CN                   C   2H   2N   1     G    300.00   3500.00 1350.00      1
 4.88864251e+00 8.97937030e-03-4.42991172e-06 1.04146368e-09-8.86722792e-14    2
 2.97135250e+04-5.23785684e-01 3.14472187e+00 1.41465426e-02-1.01712143e-05    3
 3.87667481e-09-6.13711377e-13 3.01843836e+04 8.41298194e+00                   4
CH2NH                   C   1H   3N   1     G    200.00   3500.00  700.00      1
 5.80669279e-01 1.46544725e-02-7.73860023e-06 1.97648488e-09-1.95880937e-13    2
 9.93682812e+03 1.93649675e+01 3.61447521e+00-2.68156146e-03 2.94100439e-05    3
-3.34031762e-08 1.24397123e-11 9.51209529e+03 5.81069017e+00                   4
CH3NH2                  C   1H   5N   1     G    200.00   3500.00  700.00      1
 1.20284984e-02 2.20167260e-02-1.17795639e-05 3.04373595e-09-3.04205308e-13    2
-3.36839831e+03 2.22359930e+01 3.27259113e+00 3.38493956e-03 2.81456929e-05    3
-3.49803181e-08 1.32758140e-11-3.82487708e+03 7.66862409e+00                   4
CH2NH2                  C   1H   4N   1     G    200.00   3500.00 1610.00      1
 5.12514648e+00 8.47270367e-03-2.64074253e-06 3.52691508e-10-1.53029563e-14    2
 1.56058532e+04-3.27656550e+00 1.70381411e+00 1.69729083e-02-1.05601879e-05    3
 3.63196494e-09-5.24506905e-13 1.67075222e+04 1.48587409e+01                   4
CH3NH                   C   1H   4N   1     G    200.00   3500.00  700.00      1
 1.06266683e+00 1.68343859e-02-8.55523914e-06 2.12514555e-09-2.06816967e-13    2
 2.05050909e+04 1.75854915e+01 3.52441781e+00 2.76723747e-03 2.15886504e-05    3
-2.65833207e-08 1.00462067e-11 2.01604458e+04 6.58701095e+00                   4
END
